-- generated with romgen by MikeJ
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity VIC20_KERNAL_ROM is
  port (
    CLK         : in    std_logic;
    ADDR        : in    std_logic_vector(12 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of VIC20_KERNAL_ROM is


  type ROM_ARRAY is array(0 to 8191) of std_logic_vector(7 downto 0);
  constant ROM : ROM_ARRAY := (
    x"0F",x"DC",x"A5",x"61",x"C9",x"88",x"90",x"03", -- 0x0000
    x"20",x"D4",x"DA",x"20",x"CC",x"DC",x"A5",x"07", -- 0x0008
    x"18",x"69",x"81",x"F0",x"F3",x"38",x"E9",x"01", -- 0x0010
    x"48",x"A2",x"05",x"B5",x"69",x"B4",x"61",x"95", -- 0x0018
    x"61",x"94",x"69",x"CA",x"10",x"F5",x"A5",x"56", -- 0x0020
    x"85",x"70",x"20",x"53",x"D8",x"20",x"B4",x"DF", -- 0x0028
    x"A9",x"C4",x"A0",x"DF",x"20",x"56",x"E0",x"A9", -- 0x0030
    x"00",x"85",x"6F",x"68",x"20",x"B9",x"DA",x"60", -- 0x0038
    x"85",x"71",x"84",x"72",x"20",x"CA",x"DB",x"A9", -- 0x0040
    x"57",x"20",x"28",x"DA",x"20",x"5A",x"E0",x"A9", -- 0x0048
    x"57",x"A0",x"00",x"4C",x"28",x"DA",x"85",x"71", -- 0x0050
    x"84",x"72",x"20",x"C7",x"DB",x"B1",x"71",x"85", -- 0x0058
    x"67",x"A4",x"71",x"C8",x"98",x"D0",x"02",x"E6", -- 0x0060
    x"72",x"85",x"71",x"A4",x"72",x"20",x"28",x"DA", -- 0x0068
    x"A5",x"71",x"A4",x"72",x"18",x"69",x"05",x"90", -- 0x0070
    x"01",x"C8",x"85",x"71",x"84",x"72",x"20",x"67", -- 0x0078
    x"D8",x"A9",x"5C",x"A0",x"00",x"C6",x"67",x"D0", -- 0x0080
    x"E4",x"60",x"98",x"35",x"44",x"7A",x"00",x"68", -- 0x0088
    x"28",x"B1",x"46",x"00",x"20",x"2B",x"DC",x"30", -- 0x0090
    x"37",x"D0",x"20",x"20",x"F3",x"FF",x"86",x"22", -- 0x0098
    x"84",x"23",x"A0",x"04",x"B1",x"22",x"85",x"62", -- 0x00A0
    x"C8",x"B1",x"22",x"85",x"64",x"A0",x"08",x"B1", -- 0x00A8
    x"22",x"85",x"63",x"C8",x"B1",x"22",x"85",x"65", -- 0x00B0
    x"4C",x"E0",x"E0",x"A9",x"8B",x"A0",x"00",x"20", -- 0x00B8
    x"A2",x"DB",x"A9",x"8A",x"A0",x"E0",x"20",x"28", -- 0x00C0
    x"DA",x"A9",x"8F",x"A0",x"E0",x"20",x"67",x"D8", -- 0x00C8
    x"A6",x"65",x"A5",x"62",x"85",x"65",x"86",x"62", -- 0x00D0
    x"A6",x"63",x"A5",x"64",x"85",x"63",x"86",x"64", -- 0x00D8
    x"A9",x"00",x"85",x"66",x"A5",x"61",x"85",x"70", -- 0x00E0
    x"A9",x"80",x"85",x"61",x"20",x"D7",x"D8",x"A2", -- 0x00E8
    x"8B",x"A0",x"00",x"4C",x"D4",x"DB",x"C9",x"F0", -- 0x00F0
    x"D0",x"07",x"84",x"38",x"86",x"37",x"4C",x"63", -- 0x00F8
    x"C6",x"AA",x"D0",x"02",x"A2",x"1E",x"4C",x"37", -- 0x0100
    x"C4",x"20",x"D2",x"FF",x"B0",x"E8",x"60",x"20", -- 0x0108
    x"CF",x"FF",x"B0",x"E2",x"60",x"20",x"C9",x"FF", -- 0x0110
    x"B0",x"DC",x"60",x"20",x"C6",x"FF",x"B0",x"D6", -- 0x0118
    x"60",x"20",x"E4",x"FF",x"B0",x"D0",x"60",x"20", -- 0x0120
    x"8A",x"CD",x"20",x"F7",x"D7",x"A9",x"E1",x"48", -- 0x0128
    x"A9",x"43",x"48",x"AD",x"0F",x"03",x"48",x"AD", -- 0x0130
    x"0C",x"03",x"AE",x"0D",x"03",x"AC",x"0E",x"03", -- 0x0138
    x"28",x"6C",x"14",x"00",x"08",x"8D",x"0C",x"03", -- 0x0140
    x"8E",x"0D",x"03",x"8C",x"0E",x"03",x"68",x"8D", -- 0x0148
    x"0F",x"03",x"60",x"20",x"D1",x"E1",x"A6",x"2D", -- 0x0150
    x"A4",x"2E",x"A9",x"2B",x"20",x"D8",x"FF",x"B0", -- 0x0158
    x"95",x"60",x"A9",x"01",x"2C",x"A9",x"00",x"85", -- 0x0160
    x"0A",x"20",x"D1",x"E1",x"A5",x"0A",x"A6",x"2B", -- 0x0168
    x"A4",x"2C",x"20",x"D5",x"FF",x"B0",x"57",x"A5", -- 0x0170
    x"0A",x"F0",x"1A",x"A2",x"1C",x"20",x"B7",x"FF", -- 0x0178
    x"29",x"10",x"F0",x"03",x"4C",x"37",x"C4",x"A5", -- 0x0180
    x"7A",x"C9",x"02",x"F0",x"07",x"A9",x"64",x"A0", -- 0x0188
    x"C3",x"4C",x"1E",x"CB",x"60",x"20",x"B7",x"FF", -- 0x0190
    x"29",x"BF",x"F0",x"05",x"A2",x"1D",x"4C",x"37", -- 0x0198
    x"C4",x"A5",x"7B",x"C9",x"02",x"D0",x"0E",x"86", -- 0x01A0
    x"2D",x"84",x"2E",x"A9",x"76",x"A0",x"C3",x"20", -- 0x01A8
    x"1E",x"CB",x"4C",x"2A",x"C5",x"20",x"8E",x"C6", -- 0x01B0
    x"4C",x"76",x"E4",x"20",x"16",x"E2",x"20",x"C0", -- 0x01B8
    x"FF",x"B0",x"0B",x"60",x"20",x"16",x"E2",x"A5", -- 0x01C0
    x"49",x"20",x"C3",x"FF",x"90",x"C6",x"4C",x"F6", -- 0x01C8
    x"E0",x"A9",x"00",x"20",x"BD",x"FF",x"A2",x"01", -- 0x01D0
    x"A0",x"00",x"20",x"BA",x"FF",x"20",x"03",x"E2", -- 0x01D8
    x"20",x"54",x"E2",x"20",x"03",x"E2",x"20",x"FD", -- 0x01E0
    x"E1",x"A0",x"00",x"86",x"49",x"20",x"BA",x"FF", -- 0x01E8
    x"20",x"03",x"E2",x"20",x"FD",x"E1",x"8A",x"A8", -- 0x01F0
    x"A6",x"49",x"4C",x"BA",x"FF",x"20",x"0B",x"E2", -- 0x01F8
    x"4C",x"9E",x"D7",x"20",x"79",x"00",x"D0",x"02", -- 0x0200
    x"68",x"68",x"60",x"20",x"FD",x"CE",x"20",x"79", -- 0x0208
    x"00",x"D0",x"F7",x"4C",x"08",x"CF",x"A9",x"00", -- 0x0210
    x"20",x"BD",x"FF",x"20",x"0E",x"E2",x"20",x"9E", -- 0x0218
    x"D7",x"86",x"49",x"8A",x"A2",x"01",x"A0",x"00", -- 0x0220
    x"20",x"BA",x"FF",x"20",x"03",x"E2",x"20",x"FD", -- 0x0228
    x"E1",x"86",x"4A",x"A0",x"00",x"A5",x"49",x"E0", -- 0x0230
    x"03",x"90",x"01",x"88",x"20",x"BA",x"FF",x"20", -- 0x0238
    x"03",x"E2",x"20",x"FD",x"E1",x"8A",x"A8",x"A6", -- 0x0240
    x"4A",x"A5",x"49",x"20",x"BA",x"FF",x"20",x"03", -- 0x0248
    x"E2",x"20",x"0B",x"E2",x"20",x"9E",x"CD",x"20", -- 0x0250
    x"A3",x"D6",x"A6",x"22",x"A4",x"23",x"4C",x"BD", -- 0x0258
    x"FF",x"A9",x"DD",x"A0",x"E2",x"20",x"67",x"D8", -- 0x0260
    x"20",x"0C",x"DC",x"A9",x"E2",x"A0",x"E2",x"A6", -- 0x0268
    x"6E",x"20",x"07",x"DB",x"20",x"0C",x"DC",x"20", -- 0x0270
    x"CC",x"DC",x"A9",x"00",x"85",x"6F",x"20",x"53", -- 0x0278
    x"D8",x"A9",x"E7",x"A0",x"E2",x"20",x"50",x"D8", -- 0x0280
    x"A5",x"66",x"48",x"10",x"0D",x"20",x"49",x"D8", -- 0x0288
    x"A5",x"66",x"30",x"09",x"A5",x"12",x"49",x"FF", -- 0x0290
    x"85",x"12",x"20",x"B4",x"DF",x"A9",x"E7",x"A0", -- 0x0298
    x"E2",x"20",x"67",x"D8",x"68",x"10",x"03",x"20", -- 0x02A0
    x"B4",x"DF",x"A9",x"EC",x"A0",x"E2",x"4C",x"40", -- 0x02A8
    x"E0",x"20",x"CA",x"DB",x"A9",x"00",x"85",x"12", -- 0x02B0
    x"20",x"68",x"E2",x"A2",x"4E",x"A0",x"00",x"20", -- 0x02B8
    x"F3",x"E0",x"A9",x"57",x"A0",x"00",x"20",x"A2", -- 0x02C0
    x"DB",x"A9",x"00",x"85",x"66",x"A5",x"12",x"20", -- 0x02C8
    x"D9",x"E2",x"A9",x"4E",x"A0",x"00",x"4C",x"0F", -- 0x02D0
    x"DB",x"48",x"4C",x"9A",x"E2",x"81",x"49",x"0F", -- 0x02D8
    x"DA",x"A2",x"83",x"49",x"0F",x"DA",x"A2",x"7F", -- 0x02E0
    x"00",x"00",x"00",x"00",x"05",x"84",x"E6",x"1A", -- 0x02E8
    x"2D",x"1B",x"86",x"28",x"07",x"FB",x"F8",x"87", -- 0x02F0
    x"99",x"68",x"89",x"01",x"87",x"23",x"35",x"DF", -- 0x02F8
    x"E1",x"86",x"A5",x"5D",x"E7",x"28",x"83",x"49", -- 0x0300
    x"0F",x"DA",x"A2",x"A5",x"66",x"48",x"10",x"03", -- 0x0308
    x"20",x"B4",x"DF",x"A5",x"61",x"48",x"C9",x"81", -- 0x0310
    x"90",x"07",x"A9",x"BC",x"A0",x"D9",x"20",x"0F", -- 0x0318
    x"DB",x"A9",x"3B",x"A0",x"E3",x"20",x"40",x"E0", -- 0x0320
    x"68",x"C9",x"81",x"90",x"07",x"A9",x"DD",x"A0", -- 0x0328
    x"E2",x"20",x"50",x"D8",x"68",x"10",x"03",x"4C", -- 0x0330
    x"B4",x"DF",x"60",x"0B",x"76",x"B3",x"83",x"BD", -- 0x0338
    x"D3",x"79",x"1E",x"F4",x"A6",x"F5",x"7B",x"83", -- 0x0340
    x"FC",x"B0",x"10",x"7C",x"0C",x"1F",x"67",x"CA", -- 0x0348
    x"7C",x"DE",x"53",x"CB",x"C1",x"7D",x"14",x"64", -- 0x0350
    x"70",x"4C",x"7D",x"B7",x"EA",x"51",x"7A",x"7D", -- 0x0358
    x"63",x"30",x"88",x"7E",x"7E",x"92",x"44",x"99", -- 0x0360
    x"3A",x"7E",x"4C",x"CC",x"91",x"C7",x"7F",x"AA", -- 0x0368
    x"AA",x"AA",x"13",x"81",x"00",x"00",x"00",x"00", -- 0x0370
    x"20",x"5B",x"E4",x"20",x"A4",x"E3",x"20",x"04", -- 0x0378
    x"E4",x"A2",x"FB",x"9A",x"4C",x"74",x"C4",x"E6", -- 0x0380
    x"7A",x"D0",x"02",x"E6",x"7B",x"AD",x"60",x"EA", -- 0x0388
    x"C9",x"3A",x"B0",x"0A",x"C9",x"20",x"F0",x"EF", -- 0x0390
    x"38",x"E9",x"30",x"38",x"E9",x"D0",x"60",x"80", -- 0x0398
    x"4F",x"C7",x"52",x"58",x"A9",x"4C",x"85",x"54", -- 0x03A0
    x"85",x"00",x"A9",x"48",x"A0",x"D2",x"85",x"01", -- 0x03A8
    x"84",x"02",x"A9",x"91",x"A0",x"D3",x"85",x"05", -- 0x03B0
    x"84",x"06",x"A9",x"AA",x"A0",x"D1",x"85",x"03", -- 0x03B8
    x"84",x"04",x"A2",x"1C",x"BD",x"87",x"E3",x"95", -- 0x03C0
    x"73",x"CA",x"10",x"F8",x"A9",x"03",x"85",x"53", -- 0x03C8
    x"A9",x"00",x"85",x"68",x"85",x"13",x"85",x"18", -- 0x03D0
    x"A2",x"01",x"8E",x"FD",x"01",x"8E",x"FC",x"01", -- 0x03D8
    x"A2",x"19",x"86",x"16",x"38",x"20",x"9C",x"FF", -- 0x03E0
    x"86",x"2B",x"84",x"2C",x"38",x"20",x"99",x"FF", -- 0x03E8
    x"86",x"37",x"84",x"38",x"86",x"33",x"84",x"34", -- 0x03F0
    x"A0",x"00",x"98",x"91",x"2B",x"E6",x"2B",x"D0", -- 0x03F8
    x"02",x"E6",x"2C",x"60",x"A5",x"2B",x"A4",x"2C", -- 0x0400
    x"20",x"08",x"C4",x"A9",x"36",x"A0",x"E4",x"20", -- 0x0408
    x"1E",x"CB",x"A5",x"37",x"38",x"E5",x"2B",x"AA", -- 0x0410
    x"A5",x"38",x"E5",x"2C",x"20",x"CD",x"DD",x"A9", -- 0x0418
    x"29",x"A0",x"E4",x"20",x"1E",x"CB",x"4C",x"44", -- 0x0420
    x"C6",x"20",x"42",x"59",x"54",x"45",x"53",x"20", -- 0x0428
    x"46",x"52",x"45",x"45",x"0D",x"00",x"93",x"2A", -- 0x0430
    x"2A",x"2A",x"2A",x"20",x"43",x"42",x"4D",x"20", -- 0x0438
    x"42",x"41",x"53",x"49",x"43",x"20",x"56",x"32", -- 0x0440
    x"20",x"2A",x"2A",x"2A",x"2A",x"0D",x"00",x"3A", -- 0x0448
    x"C4",x"83",x"C4",x"7C",x"C5",x"1A",x"C7",x"E4", -- 0x0450
    x"C7",x"86",x"CE",x"A2",x"0B",x"BD",x"4F",x"E4", -- 0x0458
    x"9D",x"00",x"03",x"CA",x"10",x"F7",x"60",x"20", -- 0x0460
    x"CC",x"FF",x"A9",x"00",x"85",x"13",x"20",x"7A", -- 0x0468
    x"C6",x"58",x"4C",x"74",x"C4",x"FE",x"20",x"33", -- 0x0470
    x"C5",x"4C",x"77",x"C6",x"AA",x"AA",x"AA",x"AA", -- 0x0478
    x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA", -- 0x0480
    x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA", -- 0x0488
    x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA", -- 0x0490
    x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA", -- 0x0498
    x"AD",x"2C",x"91",x"29",x"DF",x"8D",x"2C",x"91", -- 0x04A0
    x"60",x"AD",x"2C",x"91",x"09",x"20",x"8D",x"2C", -- 0x04A8
    x"91",x"60",x"AD",x"1F",x"91",x"CD",x"1F",x"91", -- 0x04B0
    x"D0",x"F8",x"4A",x"60",x"A6",x"B9",x"4C",x"47", -- 0x04B8
    x"F6",x"8A",x"D0",x"08",x"A5",x"C3",x"85",x"AE", -- 0x04C0
    x"A5",x"C4",x"85",x"AF",x"4C",x"6A",x"F6",x"AA", -- 0x04C8
    x"38",x"2E",x"20",x"91",x"AD",x"21",x"91",x"6E", -- 0x04D0
    x"20",x"91",x"29",x"40",x"F0",x"03",x"86",x"91", -- 0x04D8
    x"60",x"8A",x"29",x"FD",x"85",x"91",x"60",x"AA", -- 0x04E0
    x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA", -- 0x04E8
    x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA", -- 0x04F0
    x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA", -- 0x04F8
    x"A2",x"10",x"A0",x"91",x"60",x"A2",x"16",x"A0", -- 0x0500
    x"17",x"60",x"B0",x"07",x"86",x"D6",x"84",x"D3", -- 0x0508
    x"20",x"87",x"E5",x"A6",x"D6",x"A4",x"D3",x"60", -- 0x0510
    x"20",x"BB",x"E5",x"AD",x"88",x"02",x"29",x"FD", -- 0x0518
    x"0A",x"0A",x"09",x"80",x"8D",x"05",x"90",x"AD", -- 0x0520
    x"88",x"02",x"29",x"02",x"F0",x"08",x"A9",x"80", -- 0x0528
    x"0D",x"02",x"90",x"8D",x"02",x"90",x"A9",x"00", -- 0x0530
    x"8D",x"91",x"02",x"85",x"CF",x"A9",x"DC",x"8D", -- 0x0538
    x"8F",x"02",x"A9",x"EB",x"8D",x"90",x"02",x"A9", -- 0x0540
    x"0A",x"8D",x"89",x"02",x"8D",x"8C",x"02",x"A9", -- 0x0548
    x"06",x"8D",x"86",x"02",x"A9",x"04",x"8D",x"8B", -- 0x0550
    x"02",x"A9",x"0C",x"85",x"CD",x"85",x"CC",x"AD", -- 0x0558
    x"88",x"02",x"09",x"80",x"A8",x"A9",x"00",x"AA", -- 0x0560
    x"94",x"D9",x"18",x"69",x"16",x"90",x"01",x"C8", -- 0x0568
    x"E8",x"E0",x"18",x"D0",x"F3",x"A9",x"FF",x"95", -- 0x0570
    x"D9",x"A2",x"16",x"20",x"8D",x"EA",x"CA",x"10", -- 0x0578
    x"FA",x"A0",x"00",x"84",x"D3",x"84",x"D6",x"A6", -- 0x0580
    x"D6",x"A5",x"D3",x"B4",x"D9",x"30",x"08",x"18", -- 0x0588
    x"69",x"16",x"85",x"D3",x"CA",x"10",x"F4",x"B5", -- 0x0590
    x"D9",x"29",x"03",x"0D",x"88",x"02",x"85",x"D2", -- 0x0598
    x"BD",x"FD",x"ED",x"85",x"D1",x"A9",x"15",x"E8", -- 0x05A0
    x"B4",x"D9",x"30",x"06",x"18",x"69",x"16",x"E8", -- 0x05A8
    x"10",x"F6",x"85",x"D5",x"60",x"20",x"BB",x"E5", -- 0x05B0
    x"4C",x"81",x"E5",x"A9",x"03",x"85",x"9A",x"A9", -- 0x05B8
    x"00",x"85",x"99",x"A2",x"10",x"BD",x"E3",x"ED", -- 0x05C0
    x"9D",x"FF",x"8F",x"CA",x"D0",x"F7",x"60",x"AC", -- 0x05C8
    x"77",x"02",x"A2",x"00",x"BD",x"78",x"02",x"9D", -- 0x05D0
    x"77",x"02",x"E8",x"E4",x"C6",x"D0",x"F5",x"C6", -- 0x05D8
    x"C6",x"98",x"58",x"18",x"60",x"20",x"42",x"E7", -- 0x05E0
    x"A5",x"C6",x"85",x"CC",x"8D",x"92",x"02",x"F0", -- 0x05E8
    x"F7",x"78",x"A5",x"CF",x"F0",x"0C",x"A5",x"CE", -- 0x05F0
    x"AE",x"87",x"02",x"A0",x"00",x"84",x"CF",x"20", -- 0x05F8
    x"A1",x"EA",x"20",x"CF",x"E5",x"C9",x"83",x"D0", -- 0x0600
    x"10",x"A2",x"09",x"78",x"86",x"C6",x"BD",x"F3", -- 0x0608
    x"ED",x"9D",x"76",x"02",x"CA",x"D0",x"F7",x"F0", -- 0x0610
    x"CF",x"C9",x"0D",x"D0",x"C8",x"A4",x"D5",x"84", -- 0x0618
    x"D0",x"B1",x"D1",x"C9",x"20",x"D0",x"03",x"88", -- 0x0620
    x"D0",x"F7",x"C8",x"84",x"C8",x"A0",x"00",x"8C", -- 0x0628
    x"92",x"02",x"84",x"D3",x"84",x"D4",x"A5",x"C9", -- 0x0630
    x"30",x"1D",x"A6",x"D6",x"20",x"19",x"E7",x"E4", -- 0x0638
    x"C9",x"D0",x"14",x"D0",x"12",x"A5",x"CA",x"85", -- 0x0640
    x"D3",x"C5",x"C8",x"90",x"0A",x"B0",x"42",x"98", -- 0x0648
    x"48",x"8A",x"48",x"A5",x"D0",x"F0",x"91",x"A4", -- 0x0650
    x"D3",x"B1",x"D1",x"EA",x"EA",x"EA",x"EA",x"EA", -- 0x0658
    x"EA",x"EA",x"EA",x"EA",x"EA",x"EA",x"EA",x"EA", -- 0x0660
    x"EA",x"EA",x"EA",x"EA",x"EA",x"EA",x"EA",x"EA", -- 0x0668
    x"EA",x"EA",x"85",x"D7",x"29",x"3F",x"06",x"D7", -- 0x0670
    x"24",x"D7",x"10",x"02",x"09",x"80",x"90",x"04", -- 0x0678
    x"A6",x"D4",x"D0",x"04",x"70",x"02",x"09",x"40", -- 0x0680
    x"E6",x"D3",x"20",x"B8",x"E6",x"C4",x"C8",x"D0", -- 0x0688
    x"17",x"A9",x"00",x"85",x"D0",x"A9",x"0D",x"A6", -- 0x0690
    x"99",x"E0",x"03",x"F0",x"06",x"A6",x"9A",x"E0", -- 0x0698
    x"03",x"F0",x"03",x"20",x"42",x"E7",x"A9",x"0D", -- 0x06A0
    x"85",x"D7",x"68",x"AA",x"68",x"A8",x"A5",x"D7", -- 0x06A8
    x"C9",x"DE",x"D0",x"02",x"A9",x"FF",x"18",x"60", -- 0x06B0
    x"C9",x"22",x"D0",x"08",x"A5",x"D4",x"49",x"01", -- 0x06B8
    x"85",x"D4",x"A9",x"22",x"60",x"09",x"40",x"A6", -- 0x06C0
    x"C7",x"F0",x"02",x"09",x"80",x"A6",x"D8",x"F0", -- 0x06C8
    x"02",x"C6",x"D8",x"AE",x"86",x"02",x"20",x"A1", -- 0x06D0
    x"EA",x"20",x"EA",x"E6",x"68",x"A8",x"A5",x"D8", -- 0x06D8
    x"F0",x"02",x"46",x"D4",x"68",x"AA",x"68",x"18", -- 0x06E0
    x"58",x"60",x"20",x"FA",x"E8",x"E6",x"D3",x"A5", -- 0x06E8
    x"D5",x"C5",x"D3",x"B0",x"37",x"C9",x"57",x"F0", -- 0x06F0
    x"2A",x"AD",x"92",x"02",x"F0",x"03",x"4C",x"F0", -- 0x06F8
    x"E9",x"A6",x"D6",x"E0",x"17",x"90",x"07",x"20", -- 0x0700
    x"75",x"E9",x"C6",x"D6",x"A6",x"D6",x"16",x"D9", -- 0x0708
    x"56",x"D9",x"4C",x"5B",x"ED",x"69",x"16",x"85", -- 0x0710
    x"D5",x"B5",x"D9",x"30",x"03",x"CA",x"D0",x"F9", -- 0x0718
    x"4C",x"7E",x"EA",x"C6",x"D6",x"20",x"C3",x"E8", -- 0x0720
    x"A9",x"00",x"85",x"D3",x"60",x"A6",x"D6",x"D0", -- 0x0728
    x"06",x"86",x"D3",x"68",x"68",x"D0",x"A5",x"CA", -- 0x0730
    x"86",x"D6",x"20",x"87",x"E5",x"A4",x"D5",x"84", -- 0x0738
    x"D3",x"60",x"48",x"85",x"D7",x"8A",x"48",x"98", -- 0x0740
    x"48",x"A9",x"00",x"85",x"D0",x"A4",x"D3",x"A5", -- 0x0748
    x"D7",x"10",x"03",x"4C",x"00",x"E8",x"C9",x"0D", -- 0x0750
    x"D0",x"03",x"4C",x"D8",x"E8",x"C9",x"20",x"90", -- 0x0758
    x"10",x"C9",x"60",x"90",x"04",x"29",x"DF",x"D0", -- 0x0760
    x"02",x"29",x"3F",x"20",x"B8",x"E6",x"4C",x"C7", -- 0x0768
    x"E6",x"A6",x"D8",x"F0",x"03",x"4C",x"CB",x"E6", -- 0x0770
    x"C9",x"14",x"D0",x"2E",x"98",x"D0",x"06",x"20", -- 0x0778
    x"2D",x"E7",x"4C",x"9F",x"E7",x"20",x"E8",x"E8", -- 0x0780
    x"88",x"84",x"D3",x"20",x"B2",x"EA",x"C8",x"B1", -- 0x0788
    x"D1",x"88",x"91",x"D1",x"C8",x"B1",x"F3",x"88", -- 0x0790
    x"91",x"F3",x"C8",x"C4",x"D5",x"D0",x"EF",x"A9", -- 0x0798
    x"20",x"91",x"D1",x"AD",x"86",x"02",x"91",x"F3", -- 0x07A0
    x"10",x"4D",x"A6",x"D4",x"F0",x"03",x"4C",x"CB", -- 0x07A8
    x"E6",x"C9",x"12",x"D0",x"02",x"85",x"C7",x"C9", -- 0x07B0
    x"13",x"D0",x"03",x"20",x"81",x"E5",x"C9",x"1D", -- 0x07B8
    x"D0",x"17",x"C8",x"20",x"FA",x"E8",x"84",x"D3", -- 0x07C0
    x"88",x"C4",x"D5",x"90",x"09",x"C6",x"D6",x"20", -- 0x07C8
    x"C3",x"E8",x"A0",x"00",x"84",x"D3",x"4C",x"DC", -- 0x07D0
    x"E6",x"C9",x"11",x"D0",x"1D",x"18",x"98",x"69", -- 0x07D8
    x"16",x"A8",x"E6",x"D6",x"C5",x"D5",x"90",x"EC", -- 0x07E0
    x"F0",x"EA",x"C6",x"D6",x"E9",x"16",x"90",x"04", -- 0x07E8
    x"85",x"D3",x"D0",x"F8",x"20",x"C3",x"E8",x"4C", -- 0x07F0
    x"DC",x"E6",x"20",x"12",x"E9",x"4C",x"21",x"ED", -- 0x07F8
    x"EA",x"EA",x"EA",x"EA",x"EA",x"EA",x"EA",x"EA", -- 0x0800
    x"EA",x"EA",x"EA",x"EA",x"EA",x"EA",x"EA",x"EA", -- 0x0808
    x"EA",x"EA",x"EA",x"EA",x"EA",x"29",x"7F",x"C9", -- 0x0810
    x"7F",x"D0",x"02",x"A9",x"5E",x"EA",x"EA",x"EA", -- 0x0818
    x"EA",x"EA",x"EA",x"C9",x"20",x"90",x"03",x"4C", -- 0x0820
    x"C5",x"E6",x"C9",x"0D",x"D0",x"03",x"4C",x"D8", -- 0x0828
    x"E8",x"A6",x"D4",x"D0",x"3F",x"C9",x"14",x"D0", -- 0x0830
    x"37",x"A4",x"D5",x"B1",x"D1",x"C9",x"20",x"D0", -- 0x0838
    x"04",x"C4",x"D3",x"D0",x"07",x"C0",x"57",x"F0", -- 0x0840
    x"24",x"20",x"EE",x"E9",x"A4",x"D5",x"20",x"B2", -- 0x0848
    x"EA",x"88",x"B1",x"D1",x"C8",x"91",x"D1",x"88", -- 0x0850
    x"B1",x"F3",x"C8",x"91",x"F3",x"88",x"C4",x"D3", -- 0x0858
    x"D0",x"EF",x"A9",x"20",x"91",x"D1",x"AD",x"86", -- 0x0860
    x"02",x"91",x"F3",x"E6",x"D8",x"4C",x"DC",x"E6", -- 0x0868
    x"A6",x"D8",x"F0",x"05",x"09",x"40",x"4C",x"CB", -- 0x0870
    x"E6",x"C9",x"11",x"D0",x"16",x"A6",x"D6",x"F0", -- 0x0878
    x"37",x"C6",x"D6",x"A5",x"D3",x"38",x"E9",x"16", -- 0x0880
    x"90",x"04",x"85",x"D3",x"10",x"2A",x"20",x"87", -- 0x0888
    x"E5",x"D0",x"25",x"C9",x"12",x"D0",x"04",x"A9", -- 0x0890
    x"00",x"85",x"C7",x"C9",x"1D",x"D0",x"12",x"98", -- 0x0898
    x"F0",x"09",x"20",x"E8",x"E8",x"88",x"84",x"D3", -- 0x08A0
    x"4C",x"DC",x"E6",x"20",x"2D",x"E7",x"4C",x"DC", -- 0x08A8
    x"E6",x"C9",x"13",x"D0",x"06",x"20",x"5F",x"E5", -- 0x08B0
    x"4C",x"DC",x"E6",x"09",x"80",x"20",x"12",x"E9", -- 0x08B8
    x"4C",x"30",x"ED",x"46",x"C9",x"A6",x"D6",x"E8", -- 0x08C0
    x"E0",x"17",x"D0",x"03",x"20",x"75",x"E9",x"B5", -- 0x08C8
    x"D9",x"10",x"F4",x"86",x"D6",x"4C",x"87",x"E5", -- 0x08D0
    x"A2",x"00",x"86",x"D8",x"86",x"C7",x"86",x"D4", -- 0x08D8
    x"86",x"D3",x"20",x"C3",x"E8",x"4C",x"DC",x"E6", -- 0x08E0
    x"A2",x"04",x"A9",x"00",x"C5",x"D3",x"F0",x"07", -- 0x08E8
    x"18",x"69",x"16",x"CA",x"D0",x"F6",x"60",x"C6", -- 0x08F0
    x"D6",x"60",x"A2",x"04",x"A9",x"15",x"C5",x"D3", -- 0x08F8
    x"F0",x"07",x"18",x"69",x"16",x"CA",x"D0",x"F6", -- 0x0900
    x"60",x"A6",x"D6",x"E0",x"17",x"F0",x"02",x"E6", -- 0x0908
    x"D6",x"60",x"A2",x"07",x"DD",x"21",x"E9",x"F0", -- 0x0910
    x"04",x"CA",x"10",x"F8",x"60",x"8E",x"86",x"02", -- 0x0918
    x"60",x"90",x"05",x"1C",x"9F",x"9C",x"1E",x"1F", -- 0x0920
    x"9E",x"EF",x"A1",x"DF",x"A6",x"E1",x"B1",x"E2", -- 0x0928
    x"B2",x"E3",x"B3",x"E4",x"B4",x"E5",x"B5",x"E6", -- 0x0930
    x"B6",x"E7",x"B7",x"E8",x"B8",x"E9",x"B9",x"FA", -- 0x0938
    x"BA",x"FB",x"BB",x"FC",x"BC",x"EC",x"BD",x"FE", -- 0x0940
    x"BE",x"84",x"BF",x"F7",x"C0",x"F8",x"DB",x"F9", -- 0x0948
    x"DD",x"EA",x"DE",x"5E",x"E0",x"5B",x"E1",x"5D", -- 0x0950
    x"E2",x"40",x"B0",x"61",x"B1",x"78",x"DB",x"79", -- 0x0958
    x"DD",x"66",x"B6",x"77",x"C0",x"70",x"F0",x"71", -- 0x0960
    x"F1",x"72",x"F2",x"73",x"F3",x"74",x"F4",x"75", -- 0x0968
    x"F5",x"76",x"F6",x"7D",x"FD",x"A5",x"AC",x"48", -- 0x0970
    x"A5",x"AD",x"48",x"A5",x"AE",x"48",x"A5",x"AF", -- 0x0978
    x"48",x"A2",x"FF",x"C6",x"D6",x"C6",x"C9",x"C6", -- 0x0980
    x"F2",x"E8",x"20",x"7E",x"EA",x"E0",x"16",x"B0", -- 0x0988
    x"0C",x"BD",x"FE",x"ED",x"85",x"AC",x"B5",x"DA", -- 0x0990
    x"20",x"56",x"EA",x"30",x"EC",x"20",x"8D",x"EA", -- 0x0998
    x"A2",x"00",x"B5",x"D9",x"29",x"7F",x"B4",x"DA", -- 0x09A0
    x"10",x"02",x"09",x"80",x"95",x"D9",x"E8",x"E0", -- 0x09A8
    x"16",x"D0",x"EF",x"A5",x"EF",x"09",x"80",x"85", -- 0x09B0
    x"EF",x"A5",x"D9",x"10",x"C4",x"E6",x"D6",x"E6", -- 0x09B8
    x"F2",x"A9",x"FB",x"8D",x"20",x"91",x"AD",x"21", -- 0x09C0
    x"91",x"C9",x"FE",x"08",x"A9",x"F7",x"8D",x"20", -- 0x09C8
    x"91",x"28",x"D0",x"0B",x"A0",x"00",x"EA",x"CA", -- 0x09D0
    x"D0",x"FC",x"88",x"D0",x"F9",x"84",x"C6",x"A6", -- 0x09D8
    x"D6",x"68",x"85",x"AF",x"68",x"85",x"AE",x"68", -- 0x09E0
    x"85",x"AD",x"68",x"85",x"AC",x"60",x"A6",x"D6", -- 0x09E8
    x"E8",x"B5",x"D9",x"10",x"FB",x"86",x"F2",x"E0", -- 0x09F0
    x"16",x"F0",x"0D",x"90",x"0B",x"20",x"75",x"E9", -- 0x09F8
    x"A6",x"F2",x"CA",x"C6",x"D6",x"4C",x"0E",x"E7", -- 0x0A00
    x"A5",x"AC",x"48",x"A5",x"AD",x"48",x"A5",x"AE", -- 0x0A08
    x"48",x"A5",x"AF",x"48",x"A2",x"17",x"CA",x"20", -- 0x0A10
    x"7E",x"EA",x"E4",x"F2",x"90",x"0E",x"F0",x"0C", -- 0x0A18
    x"BD",x"FC",x"ED",x"85",x"AC",x"B5",x"D8",x"20", -- 0x0A20
    x"56",x"EA",x"30",x"EA",x"20",x"8D",x"EA",x"A2", -- 0x0A28
    x"15",x"E4",x"F2",x"90",x"0F",x"B5",x"DA",x"29", -- 0x0A30
    x"7F",x"B4",x"D9",x"10",x"02",x"09",x"80",x"95", -- 0x0A38
    x"DA",x"CA",x"D0",x"ED",x"A6",x"F2",x"20",x"0E", -- 0x0A40
    x"E7",x"68",x"85",x"AF",x"68",x"85",x"AE",x"68", -- 0x0A48
    x"85",x"AD",x"68",x"85",x"AC",x"60",x"29",x"03", -- 0x0A50
    x"0D",x"88",x"02",x"85",x"AD",x"20",x"6E",x"EA", -- 0x0A58
    x"A0",x"15",x"B1",x"AC",x"91",x"D1",x"B1",x"AE", -- 0x0A60
    x"91",x"F3",x"88",x"10",x"F5",x"60",x"20",x"B2", -- 0x0A68
    x"EA",x"A5",x"AC",x"85",x"AE",x"A5",x"AD",x"29", -- 0x0A70
    x"03",x"09",x"94",x"85",x"AF",x"60",x"BD",x"FD", -- 0x0A78
    x"ED",x"85",x"D1",x"B5",x"D9",x"29",x"03",x"0D", -- 0x0A80
    x"88",x"02",x"85",x"D2",x"60",x"A0",x"15",x"20", -- 0x0A88
    x"7E",x"EA",x"20",x"B2",x"EA",x"A9",x"20",x"91", -- 0x0A90
    x"D1",x"A9",x"01",x"91",x"F3",x"88",x"10",x"F5", -- 0x0A98
    x"60",x"A8",x"A9",x"02",x"85",x"CD",x"20",x"B2", -- 0x0AA0
    x"EA",x"98",x"A4",x"D3",x"91",x"D1",x"8A",x"91", -- 0x0AA8
    x"F3",x"60",x"A5",x"D1",x"85",x"F3",x"A5",x"D2", -- 0x0AB0
    x"29",x"03",x"09",x"94",x"85",x"F4",x"60",x"20", -- 0x0AB8
    x"EA",x"FF",x"A5",x"CC",x"D0",x"29",x"C6",x"CD", -- 0x0AC0
    x"D0",x"25",x"A9",x"14",x"85",x"CD",x"A4",x"D3", -- 0x0AC8
    x"46",x"CF",x"AE",x"87",x"02",x"B1",x"D1",x"B0", -- 0x0AD0
    x"11",x"E6",x"CF",x"85",x"CE",x"20",x"B2",x"EA", -- 0x0AD8
    x"B1",x"F3",x"8D",x"87",x"02",x"AE",x"86",x"02", -- 0x0AE0
    x"A5",x"CE",x"49",x"80",x"20",x"AA",x"EA",x"AD", -- 0x0AE8
    x"1F",x"91",x"29",x"40",x"F0",x"0B",x"A0",x"00", -- 0x0AF0
    x"84",x"C0",x"AD",x"1C",x"91",x"09",x"02",x"D0", -- 0x0AF8
    x"09",x"A5",x"C0",x"D0",x"0D",x"AD",x"1C",x"91", -- 0x0B00
    x"29",x"FD",x"2C",x"1E",x"91",x"70",x"03",x"8D", -- 0x0B08
    x"1C",x"91",x"20",x"1E",x"EB",x"2C",x"24",x"91", -- 0x0B10
    x"68",x"A8",x"68",x"AA",x"68",x"40",x"A9",x"00", -- 0x0B18
    x"8D",x"8D",x"02",x"A0",x"40",x"84",x"CB",x"8D", -- 0x0B20
    x"20",x"91",x"AE",x"21",x"91",x"E0",x"FF",x"F0", -- 0x0B28
    x"5E",x"A9",x"FE",x"8D",x"20",x"91",x"A0",x"00", -- 0x0B30
    x"A9",x"5E",x"85",x"F5",x"A9",x"EC",x"85",x"F6", -- 0x0B38
    x"A2",x"08",x"AD",x"21",x"91",x"CD",x"21",x"91", -- 0x0B40
    x"D0",x"F6",x"4A",x"B0",x"16",x"48",x"B1",x"F5", -- 0x0B48
    x"C9",x"05",x"B0",x"0C",x"C9",x"03",x"F0",x"08", -- 0x0B50
    x"0D",x"8D",x"02",x"8D",x"8D",x"02",x"10",x"02", -- 0x0B58
    x"84",x"CB",x"68",x"C8",x"C0",x"41",x"B0",x"09", -- 0x0B60
    x"CA",x"D0",x"DF",x"38",x"2E",x"20",x"91",x"D0", -- 0x0B68
    x"CF",x"6C",x"8F",x"02",x"A4",x"CB",x"B1",x"F5", -- 0x0B70
    x"AA",x"C4",x"C5",x"F0",x"07",x"A0",x"10",x"8C", -- 0x0B78
    x"8C",x"02",x"D0",x"36",x"29",x"7F",x"2C",x"8A", -- 0x0B80
    x"02",x"30",x"16",x"70",x"49",x"C9",x"7F",x"F0", -- 0x0B88
    x"29",x"C9",x"14",x"F0",x"0C",x"C9",x"20",x"F0", -- 0x0B90
    x"08",x"C9",x"1D",x"F0",x"04",x"C9",x"11",x"D0", -- 0x0B98
    x"35",x"AC",x"8C",x"02",x"F0",x"05",x"CE",x"8C", -- 0x0BA0
    x"02",x"D0",x"2B",x"CE",x"8B",x"02",x"D0",x"26", -- 0x0BA8
    x"A0",x"04",x"8C",x"8B",x"02",x"A4",x"C6",x"88", -- 0x0BB0
    x"10",x"1C",x"A4",x"CB",x"84",x"C5",x"AC",x"8D", -- 0x0BB8
    x"02",x"8C",x"8E",x"02",x"E0",x"FF",x"F0",x"0E", -- 0x0BC0
    x"8A",x"A6",x"C6",x"EC",x"89",x"02",x"B0",x"06", -- 0x0BC8
    x"9D",x"77",x"02",x"E8",x"86",x"C6",x"A9",x"F7", -- 0x0BD0
    x"8D",x"20",x"91",x"60",x"AD",x"8D",x"02",x"C9", -- 0x0BD8
    x"03",x"D0",x"2C",x"CD",x"8E",x"02",x"F0",x"EE", -- 0x0BE0
    x"AD",x"91",x"02",x"30",x"56",x"EA",x"EA",x"EA", -- 0x0BE8
    x"EA",x"EA",x"EA",x"EA",x"EA",x"EA",x"EA",x"EA", -- 0x0BF0
    x"EA",x"EA",x"EA",x"EA",x"EA",x"EA",x"EA",x"EA", -- 0x0BF8
    x"AD",x"05",x"90",x"49",x"02",x"8D",x"05",x"90", -- 0x0C00
    x"EA",x"EA",x"EA",x"EA",x"4C",x"43",x"EC",x"0A", -- 0x0C08
    x"C9",x"08",x"90",x"04",x"A9",x"06",x"EA",x"EA", -- 0x0C10
    x"EA",x"EA",x"EA",x"EA",x"EA",x"EA",x"EA",x"EA", -- 0x0C18
    x"EA",x"EA",x"EA",x"EA",x"EA",x"EA",x"EA",x"EA", -- 0x0C20
    x"EA",x"EA",x"EA",x"EA",x"EA",x"EA",x"EA",x"EA", -- 0x0C28
    x"EA",x"EA",x"EA",x"EA",x"EA",x"EA",x"EA",x"EA", -- 0x0C30
    x"AA",x"BD",x"46",x"EC",x"85",x"F5",x"BD",x"47", -- 0x0C38
    x"EC",x"85",x"F6",x"4C",x"74",x"EB",x"5E",x"EC", -- 0x0C40
    x"9F",x"EC",x"E0",x"EC",x"A3",x"ED",x"5E",x"EC", -- 0x0C48
    x"9F",x"EC",x"69",x"ED",x"A3",x"ED",x"21",x"ED", -- 0x0C50
    x"69",x"ED",x"69",x"ED",x"A3",x"ED",x"31",x"33", -- 0x0C58
    x"35",x"37",x"39",x"2D",x"3A",x"14",x"5F",x"57", -- 0x0C60
    x"52",x"59",x"49",x"50",x"40",x"0D",x"04",x"41", -- 0x0C68
    x"44",x"47",x"4A",x"4C",x"5B",x"1D",x"03",x"01", -- 0x0C70
    x"58",x"56",x"4E",x"2C",x"2F",x"11",x"20",x"5A", -- 0x0C78
    x"43",x"42",x"4D",x"2E",x"01",x"85",x"02",x"53", -- 0x0C80
    x"46",x"48",x"4B",x"5C",x"3B",x"86",x"51",x"45", -- 0x0C88
    x"54",x"55",x"4F",x"5D",x"5E",x"87",x"32",x"34", -- 0x0C90
    x"36",x"38",x"30",x"3D",x"13",x"88",x"FF",x"21", -- 0x0C98
    x"23",x"25",x"27",x"29",x"C0",x"2A",x"94",x"5F", -- 0x0CA0
    x"D7",x"D2",x"D9",x"C9",x"D0",x"BA",x"8D",x"04", -- 0x0CA8
    x"C1",x"C4",x"C7",x"CA",x"CC",x"DB",x"9D",x"83", -- 0x0CB0
    x"01",x"D8",x"D6",x"CE",x"3C",x"3F",x"91",x"A0", -- 0x0CB8
    x"DA",x"C3",x"C2",x"CD",x"3E",x"01",x"89",x"02", -- 0x0CC0
    x"D3",x"C6",x"C8",x"CB",x"DC",x"2B",x"8A",x"D1", -- 0x0CC8
    x"C5",x"D4",x"D5",x"CF",x"DD",x"DE",x"8B",x"22", -- 0x0CD0
    x"24",x"26",x"28",x"30",x"3D",x"93",x"8C",x"FF", -- 0x0CD8
    x"21",x"23",x"25",x"27",x"29",x"DF",x"2A",x"94", -- 0x0CE0
    x"5F",x"B3",x"B2",x"B7",x"A2",x"AF",x"A4",x"8D", -- 0x0CE8
    x"04",x"B0",x"AC",x"A5",x"B5",x"B6",x"A8",x"9D", -- 0x0CF0
    x"83",x"01",x"BD",x"BE",x"AA",x"3C",x"3F",x"91", -- 0x0CF8
    x"A0",x"AD",x"BC",x"BF",x"A7",x"3E",x"01",x"89", -- 0x0D00
    x"02",x"AE",x"BB",x"B4",x"A1",x"A9",x"2B",x"8A", -- 0x0D08
    x"AB",x"B1",x"A3",x"B8",x"B9",x"A6",x"DE",x"8B", -- 0x0D10
    x"22",x"24",x"26",x"28",x"30",x"3D",x"93",x"8C", -- 0x0D18
    x"FF",x"C9",x"0E",x"D0",x"0B",x"A9",x"02",x"0D", -- 0x0D20
    x"05",x"90",x"8D",x"05",x"90",x"4C",x"DC",x"E6", -- 0x0D28
    x"C9",x"8E",x"D0",x"0B",x"A9",x"FD",x"2D",x"05", -- 0x0D30
    x"90",x"8D",x"05",x"90",x"4C",x"DC",x"E6",x"C9", -- 0x0D38
    x"08",x"D0",x"0A",x"A9",x"80",x"0D",x"91",x"02", -- 0x0D40
    x"8D",x"91",x"02",x"30",x"EF",x"C9",x"09",x"D0", -- 0x0D48
    x"EB",x"A9",x"7F",x"2D",x"91",x"02",x"8D",x"91", -- 0x0D50
    x"02",x"10",x"E1",x"E8",x"B5",x"D9",x"09",x"80", -- 0x0D58
    x"95",x"D9",x"CA",x"A5",x"D5",x"18",x"4C",x"15", -- 0x0D60
    x"E7",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA", -- 0x0D68
    x"AA",x"AA",x"04",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0D70
    x"E2",x"9D",x"83",x"01",x"FF",x"FF",x"FF",x"FF", -- 0x0D78
    x"FF",x"91",x"A0",x"FF",x"FF",x"FF",x"FF",x"EE", -- 0x0D80
    x"01",x"89",x"02",x"FF",x"FF",x"FF",x"FF",x"E1", -- 0x0D88
    x"FD",x"8A",x"FF",x"FF",x"FF",x"FF",x"FF",x"B0", -- 0x0D90
    x"E0",x"8B",x"F2",x"F4",x"F6",x"FF",x"F0",x"ED", -- 0x0D98
    x"93",x"8C",x"FF",x"90",x"1C",x"9C",x"1F",x"12", -- 0x0DA0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"12",x"FF",x"FF", -- 0x0DA8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0DB0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0DB8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0DC0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0DC8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0DD0
    x"FF",x"FF",x"FF",x"05",x"9F",x"1E",x"9E",x"92", -- 0x0DD8
    x"FF",x"FF",x"FF",x"FF",x"0C",x"26",x"16",x"2E", -- 0x0DE0
    x"00",x"C0",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0DE8
    x"00",x"00",x"00",x"1B",x"4C",x"4F",x"41",x"44", -- 0x0DF0
    x"0D",x"52",x"55",x"4E",x"0D",x"00",x"16",x"2C", -- 0x0DF8
    x"42",x"58",x"6E",x"84",x"9A",x"B0",x"C6",x"DC", -- 0x0E00
    x"F2",x"08",x"1E",x"34",x"4A",x"60",x"76",x"8C", -- 0x0E08
    x"A2",x"B8",x"CE",x"E4",x"09",x"40",x"2C",x"09", -- 0x0E10
    x"20",x"20",x"60",x"F1",x"48",x"24",x"94",x"10", -- 0x0E18
    x"0A",x"38",x"66",x"A3",x"20",x"49",x"EE",x"46", -- 0x0E20
    x"94",x"46",x"A3",x"68",x"85",x"95",x"20",x"A0", -- 0x0E28
    x"E4",x"C9",x"3F",x"D0",x"03",x"20",x"84",x"EF", -- 0x0E30
    x"AD",x"1F",x"91",x"09",x"80",x"8D",x"1F",x"91", -- 0x0E38
    x"20",x"8D",x"EF",x"20",x"A0",x"E4",x"20",x"96", -- 0x0E40
    x"EF",x"78",x"20",x"A0",x"E4",x"20",x"B2",x"E4", -- 0x0E48
    x"4A",x"B0",x"61",x"20",x"84",x"EF",x"24",x"A3", -- 0x0E50
    x"10",x"0C",x"20",x"B2",x"E4",x"4A",x"90",x"FA", -- 0x0E58
    x"20",x"B2",x"E4",x"4A",x"B0",x"FA",x"20",x"B2", -- 0x0E60
    x"E4",x"4A",x"90",x"FA",x"20",x"8D",x"EF",x"A9", -- 0x0E68
    x"08",x"85",x"A5",x"AD",x"1F",x"91",x"CD",x"1F", -- 0x0E70
    x"91",x"D0",x"F8",x"4A",x"4A",x"90",x"38",x"66", -- 0x0E78
    x"95",x"B0",x"05",x"20",x"A9",x"E4",x"D0",x"03", -- 0x0E80
    x"20",x"A0",x"E4",x"20",x"84",x"EF",x"EA",x"EA", -- 0x0E88
    x"EA",x"EA",x"AD",x"2C",x"91",x"29",x"DF",x"09", -- 0x0E90
    x"02",x"8D",x"2C",x"91",x"C6",x"A5",x"D0",x"D3", -- 0x0E98
    x"A9",x"04",x"8D",x"29",x"91",x"AD",x"2D",x"91", -- 0x0EA0
    x"29",x"20",x"D0",x"0B",x"20",x"B2",x"E4",x"4A", -- 0x0EA8
    x"B0",x"F3",x"58",x"60",x"A9",x"80",x"2C",x"A9", -- 0x0EB0
    x"03",x"20",x"6A",x"FE",x"58",x"18",x"90",x"49", -- 0x0EB8
    x"85",x"95",x"20",x"40",x"EE",x"AD",x"1F",x"91", -- 0x0EC0
    x"29",x"7F",x"8D",x"1F",x"91",x"60",x"85",x"95", -- 0x0EC8
    x"20",x"40",x"EE",x"78",x"20",x"A9",x"E4",x"20", -- 0x0ED0
    x"C5",x"EE",x"20",x"84",x"EF",x"20",x"B2",x"E4", -- 0x0ED8
    x"B0",x"FB",x"58",x"60",x"24",x"94",x"30",x"05", -- 0x0EE0
    x"38",x"66",x"94",x"D0",x"05",x"48",x"20",x"49", -- 0x0EE8
    x"EE",x"68",x"85",x"95",x"18",x"60",x"20",x"8D", -- 0x0EF0
    x"EF",x"AD",x"1F",x"91",x"09",x"80",x"8D",x"1F", -- 0x0EF8
    x"91",x"A9",x"5F",x"2C",x"A9",x"3F",x"20",x"1C", -- 0x0F00
    x"EE",x"20",x"C5",x"EE",x"8A",x"A2",x"0B",x"CA", -- 0x0F08
    x"D0",x"FD",x"AA",x"20",x"84",x"EF",x"4C",x"A0", -- 0x0F10
    x"E4",x"78",x"A9",x"00",x"85",x"A5",x"20",x"84", -- 0x0F18
    x"EF",x"20",x"B2",x"E4",x"90",x"FB",x"20",x"A0", -- 0x0F20
    x"E4",x"A9",x"01",x"8D",x"29",x"91",x"AD",x"2D", -- 0x0F28
    x"91",x"29",x"20",x"D0",x"07",x"20",x"B2",x"E4", -- 0x0F30
    x"B0",x"F4",x"90",x"18",x"A5",x"A5",x"F0",x"05", -- 0x0F38
    x"A9",x"02",x"4C",x"B9",x"EE",x"20",x"A9",x"E4", -- 0x0F40
    x"20",x"0C",x"EF",x"A9",x"40",x"20",x"6A",x"FE", -- 0x0F48
    x"E6",x"A5",x"D0",x"D5",x"A9",x"08",x"85",x"A5", -- 0x0F50
    x"AD",x"1F",x"91",x"CD",x"1F",x"91",x"D0",x"F8", -- 0x0F58
    x"4A",x"90",x"F5",x"4A",x"66",x"A4",x"AD",x"1F", -- 0x0F60
    x"91",x"CD",x"1F",x"91",x"D0",x"F8",x"4A",x"B0", -- 0x0F68
    x"F5",x"C6",x"A5",x"D0",x"E3",x"20",x"A9",x"E4", -- 0x0F70
    x"A5",x"90",x"F0",x"03",x"20",x"0C",x"EF",x"A5", -- 0x0F78
    x"A4",x"58",x"18",x"60",x"AD",x"2C",x"91",x"29", -- 0x0F80
    x"FD",x"8D",x"2C",x"91",x"60",x"AD",x"2C",x"91", -- 0x0F88
    x"09",x"02",x"8D",x"2C",x"91",x"60",x"A9",x"04", -- 0x0F90
    x"8D",x"29",x"91",x"AD",x"2D",x"91",x"29",x"20", -- 0x0F98
    x"F0",x"F9",x"60",x"A5",x"B4",x"F0",x"47",x"30", -- 0x0FA0
    x"3F",x"46",x"B6",x"A2",x"00",x"90",x"01",x"CA", -- 0x0FA8
    x"8A",x"45",x"BD",x"85",x"BD",x"C6",x"B4",x"F0", -- 0x0FB0
    x"06",x"8A",x"29",x"20",x"85",x"B5",x"60",x"A9", -- 0x0FB8
    x"20",x"2C",x"94",x"02",x"F0",x"14",x"30",x"1C", -- 0x0FC0
    x"70",x"14",x"A5",x"BD",x"D0",x"01",x"CA",x"C6", -- 0x0FC8
    x"B4",x"AD",x"93",x"02",x"10",x"E3",x"C6",x"B4", -- 0x0FD0
    x"D0",x"DF",x"E6",x"B4",x"D0",x"F0",x"A5",x"BD", -- 0x0FD8
    x"F0",x"ED",x"D0",x"EA",x"70",x"E9",x"50",x"E6", -- 0x0FE0
    x"E6",x"B4",x"A2",x"FF",x"D0",x"CB",x"AD",x"94", -- 0x0FE8
    x"02",x"4A",x"90",x"07",x"2C",x"20",x"91",x"10", -- 0x0FF0
    x"1D",x"50",x"1E",x"A9",x"00",x"85",x"BD",x"85", -- 0x0FF8
    x"B5",x"AE",x"98",x"02",x"86",x"B4",x"AC",x"9D", -- 0x1000
    x"02",x"CC",x"9E",x"02",x"F0",x"13",x"B1",x"F9", -- 0x1008
    x"85",x"B6",x"EE",x"9D",x"02",x"60",x"A9",x"40", -- 0x1010
    x"2C",x"A9",x"10",x"0D",x"97",x"02",x"8D",x"97", -- 0x1018
    x"02",x"A9",x"40",x"8D",x"1E",x"91",x"60",x"A2", -- 0x1020
    x"09",x"A9",x"20",x"2C",x"93",x"02",x"F0",x"01", -- 0x1028
    x"CA",x"50",x"02",x"CA",x"CA",x"60",x"A6",x"A9", -- 0x1030
    x"D0",x"2E",x"C6",x"A8",x"F0",x"31",x"30",x"0D", -- 0x1038
    x"A5",x"A7",x"45",x"AB",x"85",x"AB",x"46",x"A7", -- 0x1040
    x"66",x"AA",x"60",x"C6",x"A8",x"A5",x"A7",x"F0", -- 0x1048
    x"62",x"AD",x"93",x"02",x"0A",x"A9",x"01",x"65", -- 0x1050
    x"A8",x"D0",x"EF",x"A9",x"90",x"8D",x"1E",x"91", -- 0x1058
    x"85",x"A9",x"A9",x"20",x"8D",x"1E",x"91",x"60", -- 0x1060
    x"A5",x"A7",x"D0",x"EF",x"85",x"A9",x"60",x"AC", -- 0x1068
    x"9B",x"02",x"C8",x"CC",x"9C",x"02",x"F0",x"2A", -- 0x1070
    x"8C",x"9B",x"02",x"88",x"A5",x"AA",x"AE",x"98", -- 0x1078
    x"02",x"E0",x"09",x"F0",x"04",x"4A",x"E8",x"D0", -- 0x1080
    x"F8",x"91",x"F7",x"A9",x"20",x"2C",x"94",x"02", -- 0x1088
    x"F0",x"B9",x"30",x"B6",x"A5",x"A7",x"45",x"AB", -- 0x1090
    x"F0",x"03",x"70",x"AE",x"2C",x"50",x"AB",x"A9", -- 0x1098
    x"01",x"2C",x"A9",x"04",x"2C",x"A9",x"80",x"2C", -- 0x10A0
    x"A9",x"02",x"0D",x"97",x"02",x"8D",x"97",x"02", -- 0x10A8
    x"4C",x"5B",x"F0",x"A5",x"AA",x"D0",x"F1",x"F0", -- 0x10B0
    x"EC",x"4C",x"96",x"F7",x"85",x"9A",x"AD",x"94", -- 0x10B8
    x"02",x"4A",x"90",x"27",x"A9",x"02",x"2C",x"10", -- 0x10C0
    x"91",x"10",x"1D",x"D0",x"1E",x"AD",x"1E",x"91", -- 0x10C8
    x"29",x"30",x"D0",x"F9",x"2C",x"10",x"91",x"70", -- 0x10D0
    x"FB",x"AD",x"10",x"91",x"09",x"02",x"8D",x"10", -- 0x10D8
    x"91",x"2C",x"10",x"91",x"70",x"05",x"30",x"F9", -- 0x10E0
    x"20",x"16",x"F0",x"18",x"60",x"AC",x"9E",x"02", -- 0x10E8
    x"C8",x"CC",x"9D",x"02",x"F0",x"F7",x"8C",x"9E", -- 0x10F0
    x"02",x"88",x"91",x"F9",x"2C",x"1E",x"91",x"50", -- 0x10F8
    x"01",x"60",x"AD",x"99",x"02",x"8D",x"14",x"91", -- 0x1100
    x"AD",x"9A",x"02",x"8D",x"15",x"91",x"A9",x"C0", -- 0x1108
    x"8D",x"1E",x"91",x"4C",x"EE",x"EF",x"85",x"99", -- 0x1110
    x"AD",x"94",x"02",x"4A",x"90",x"28",x"29",x"08", -- 0x1118
    x"F0",x"24",x"A9",x"02",x"2C",x"10",x"91",x"10", -- 0x1120
    x"BF",x"F0",x"19",x"2C",x"1E",x"91",x"70",x"FB", -- 0x1128
    x"AD",x"10",x"91",x"29",x"FD",x"8D",x"10",x"91", -- 0x1130
    x"AD",x"10",x"91",x"29",x"04",x"F0",x"F9",x"A9", -- 0x1138
    x"90",x"8D",x"1E",x"91",x"18",x"60",x"AD",x"1E", -- 0x1140
    x"91",x"29",x"30",x"F0",x"F2",x"18",x"60",x"AC", -- 0x1148
    x"9C",x"02",x"CC",x"9B",x"02",x"F0",x"06",x"B1", -- 0x1150
    x"F7",x"EE",x"9C",x"02",x"60",x"A9",x"00",x"60", -- 0x1158
    x"48",x"AD",x"1E",x"91",x"F0",x"0C",x"AD",x"1E", -- 0x1160
    x"91",x"29",x"60",x"D0",x"F9",x"A9",x"10",x"8D", -- 0x1168
    x"1E",x"91",x"68",x"60",x"0D",x"49",x"2F",x"4F", -- 0x1170
    x"20",x"45",x"52",x"52",x"4F",x"52",x"20",x"A3", -- 0x1178
    x"0D",x"53",x"45",x"41",x"52",x"43",x"48",x"49", -- 0x1180
    x"4E",x"47",x"A0",x"46",x"4F",x"52",x"A0",x"0D", -- 0x1188
    x"50",x"52",x"45",x"53",x"53",x"20",x"50",x"4C", -- 0x1190
    x"41",x"59",x"20",x"4F",x"4E",x"20",x"54",x"41", -- 0x1198
    x"50",x"C5",x"50",x"52",x"45",x"53",x"53",x"20", -- 0x11A0
    x"52",x"45",x"43",x"4F",x"52",x"44",x"20",x"26", -- 0x11A8
    x"20",x"50",x"4C",x"41",x"59",x"20",x"4F",x"4E", -- 0x11B0
    x"20",x"54",x"41",x"50",x"C5",x"0D",x"4C",x"4F", -- 0x11B8
    x"41",x"44",x"49",x"4E",x"C7",x"0D",x"53",x"41", -- 0x11C0
    x"56",x"49",x"4E",x"47",x"A0",x"0D",x"56",x"45", -- 0x11C8
    x"52",x"49",x"46",x"59",x"49",x"4E",x"C7",x"0D", -- 0x11D0
    x"46",x"4F",x"55",x"4E",x"44",x"A0",x"0D",x"4F", -- 0x11D8
    x"4B",x"8D",x"24",x"9D",x"10",x"0D",x"B9",x"74", -- 0x11E0
    x"F1",x"08",x"29",x"7F",x"20",x"D2",x"FF",x"C8", -- 0x11E8
    x"28",x"10",x"F3",x"18",x"60",x"A5",x"99",x"D0", -- 0x11F0
    x"08",x"A5",x"C6",x"F0",x"6D",x"78",x"4C",x"CF", -- 0x11F8
    x"E5",x"C9",x"02",x"D0",x"18",x"84",x"97",x"20", -- 0x1200
    x"4F",x"F1",x"A4",x"97",x"18",x"60",x"A5",x"99", -- 0x1208
    x"D0",x"0B",x"A5",x"D3",x"85",x"CA",x"A5",x"D6", -- 0x1210
    x"85",x"C9",x"4C",x"4F",x"E6",x"C9",x"03",x"D0", -- 0x1218
    x"09",x"85",x"D0",x"A5",x"D5",x"85",x"C8",x"4C", -- 0x1220
    x"4F",x"E6",x"B0",x"38",x"C9",x"02",x"F0",x"3F", -- 0x1228
    x"86",x"97",x"20",x"50",x"F2",x"B0",x"16",x"48", -- 0x1230
    x"20",x"50",x"F2",x"B0",x"0D",x"D0",x"05",x"A9", -- 0x1238
    x"40",x"20",x"6A",x"FE",x"C6",x"A6",x"A6",x"97", -- 0x1240
    x"68",x"60",x"AA",x"68",x"8A",x"A6",x"97",x"60", -- 0x1248
    x"20",x"8A",x"F8",x"D0",x"0B",x"20",x"C0",x"F8", -- 0x1250
    x"B0",x"11",x"A9",x"00",x"85",x"A6",x"F0",x"F0", -- 0x1258
    x"B1",x"B2",x"18",x"60",x"A5",x"90",x"F0",x"04", -- 0x1260
    x"A9",x"0D",x"18",x"60",x"4C",x"19",x"EF",x"20", -- 0x1268
    x"05",x"F2",x"B0",x"05",x"C9",x"00",x"F0",x"F7", -- 0x1270
    x"18",x"60",x"48",x"A5",x"9A",x"C9",x"03",x"D0", -- 0x1278
    x"04",x"68",x"4C",x"42",x"E7",x"90",x"04",x"68", -- 0x1280
    x"4C",x"E4",x"EE",x"C9",x"02",x"F0",x"2A",x"68", -- 0x1288
    x"85",x"9E",x"48",x"8A",x"48",x"98",x"48",x"20", -- 0x1290
    x"8A",x"F8",x"D0",x"0E",x"20",x"E3",x"F8",x"B0", -- 0x1298
    x"0E",x"A9",x"02",x"A0",x"00",x"91",x"B2",x"C8", -- 0x12A0
    x"84",x"A6",x"A5",x"9E",x"91",x"B2",x"18",x"68", -- 0x12A8
    x"A8",x"68",x"AA",x"68",x"90",x"02",x"A9",x"00", -- 0x12B0
    x"60",x"68",x"86",x"97",x"84",x"9E",x"20",x"ED", -- 0x12B8
    x"F0",x"A6",x"97",x"A4",x"9E",x"18",x"60",x"20", -- 0x12C0
    x"CF",x"F3",x"F0",x"03",x"4C",x"84",x"F7",x"20", -- 0x12C8
    x"DF",x"F3",x"A5",x"BA",x"F0",x"16",x"C9",x"03", -- 0x12D0
    x"F0",x"12",x"B0",x"14",x"C9",x"02",x"D0",x"03", -- 0x12D8
    x"4C",x"16",x"F1",x"A6",x"B9",x"E0",x"60",x"F0", -- 0x12E0
    x"03",x"4C",x"8D",x"F7",x"85",x"99",x"18",x"60", -- 0x12E8
    x"AA",x"20",x"14",x"EE",x"A5",x"B9",x"10",x"06", -- 0x12F0
    x"20",x"D3",x"EE",x"4C",x"01",x"F3",x"20",x"CE", -- 0x12F8
    x"EE",x"8A",x"24",x"90",x"10",x"E6",x"4C",x"8A", -- 0x1300
    x"F7",x"20",x"CF",x"F3",x"F0",x"03",x"4C",x"84", -- 0x1308
    x"F7",x"20",x"DF",x"F3",x"A5",x"BA",x"D0",x"03", -- 0x1310
    x"4C",x"90",x"F7",x"C9",x"03",x"F0",x"0F",x"B0", -- 0x1318
    x"11",x"C9",x"02",x"D0",x"03",x"4C",x"BC",x"F0", -- 0x1320
    x"A6",x"B9",x"E0",x"60",x"F0",x"EA",x"85",x"9A", -- 0x1328
    x"18",x"60",x"AA",x"20",x"17",x"EE",x"A5",x"B9", -- 0x1330
    x"10",x"05",x"20",x"C5",x"EE",x"D0",x"03",x"20", -- 0x1338
    x"C0",x"EE",x"8A",x"24",x"90",x"10",x"E7",x"4C", -- 0x1340
    x"8A",x"F7",x"20",x"D4",x"F3",x"F0",x"02",x"18", -- 0x1348
    x"60",x"20",x"DF",x"F3",x"8A",x"48",x"A5",x"BA", -- 0x1350
    x"F0",x"57",x"C9",x"03",x"F0",x"53",x"B0",x"4E", -- 0x1358
    x"C9",x"02",x"D0",x"29",x"68",x"20",x"B2",x"F3", -- 0x1360
    x"A9",x"7D",x"8D",x"1E",x"91",x"A9",x"06",x"8D", -- 0x1368
    x"10",x"91",x"A9",x"EE",x"8D",x"1C",x"91",x"20", -- 0x1370
    x"75",x"FE",x"A5",x"F8",x"F0",x"01",x"C8",x"A5", -- 0x1378
    x"FA",x"F0",x"01",x"C8",x"A9",x"00",x"85",x"F8", -- 0x1380
    x"85",x"FA",x"4C",x"3C",x"F5",x"A5",x"B9",x"29", -- 0x1388
    x"0F",x"F0",x"1E",x"20",x"4D",x"F8",x"A9",x"00", -- 0x1390
    x"20",x"90",x"F2",x"4C",x"CF",x"E4",x"B0",x"2E", -- 0x1398
    x"A5",x"B9",x"C9",x"62",x"D0",x"0B",x"A9",x"05", -- 0x13A0
    x"20",x"E7",x"F7",x"4C",x"B1",x"F3",x"20",x"DA", -- 0x13A8
    x"F6",x"68",x"AA",x"C6",x"98",x"E4",x"98",x"F0", -- 0x13B0
    x"14",x"A4",x"98",x"B9",x"59",x"02",x"9D",x"59", -- 0x13B8
    x"02",x"B9",x"63",x"02",x"9D",x"63",x"02",x"B9", -- 0x13C0
    x"6D",x"02",x"9D",x"6D",x"02",x"18",x"60",x"A9", -- 0x13C8
    x"00",x"85",x"90",x"8A",x"A6",x"98",x"CA",x"30", -- 0x13D0
    x"15",x"DD",x"59",x"02",x"D0",x"F8",x"60",x"BD", -- 0x13D8
    x"59",x"02",x"85",x"B8",x"BD",x"63",x"02",x"85", -- 0x13E0
    x"BA",x"BD",x"6D",x"02",x"85",x"B9",x"60",x"A9", -- 0x13E8
    x"00",x"85",x"98",x"A2",x"03",x"E4",x"9A",x"B0", -- 0x13F0
    x"03",x"20",x"04",x"EF",x"E4",x"99",x"B0",x"03", -- 0x13F8
    x"20",x"F6",x"EE",x"86",x"9A",x"A9",x"00",x"85", -- 0x1400
    x"99",x"60",x"A6",x"B8",x"D0",x"03",x"4C",x"8D", -- 0x1408
    x"F7",x"20",x"CF",x"F3",x"D0",x"03",x"4C",x"81", -- 0x1410
    x"F7",x"A6",x"98",x"E0",x"0A",x"90",x"03",x"4C", -- 0x1418
    x"7E",x"F7",x"E6",x"98",x"A5",x"B8",x"9D",x"59", -- 0x1420
    x"02",x"A5",x"B9",x"09",x"60",x"85",x"B9",x"9D", -- 0x1428
    x"6D",x"02",x"A5",x"BA",x"9D",x"63",x"02",x"F0", -- 0x1430
    x"5A",x"C9",x"03",x"F0",x"56",x"90",x"05",x"20", -- 0x1438
    x"95",x"F4",x"90",x"4F",x"C9",x"02",x"D0",x"03", -- 0x1440
    x"4C",x"C7",x"F4",x"20",x"4D",x"F8",x"B0",x"03", -- 0x1448
    x"4C",x"96",x"F7",x"A5",x"B9",x"29",x"0F",x"D0", -- 0x1450
    x"1F",x"20",x"94",x"F8",x"B0",x"36",x"20",x"47", -- 0x1458
    x"F6",x"A5",x"B7",x"F0",x"0A",x"20",x"67",x"F8", -- 0x1460
    x"90",x"18",x"F0",x"28",x"4C",x"87",x"F7",x"20", -- 0x1468
    x"AF",x"F7",x"F0",x"20",x"90",x"0C",x"B0",x"F4", -- 0x1470
    x"20",x"B7",x"F8",x"B0",x"17",x"A9",x"04",x"20", -- 0x1478
    x"E7",x"F7",x"A9",x"BF",x"A4",x"B9",x"C0",x"60", -- 0x1480
    x"F0",x"07",x"A0",x"00",x"A9",x"02",x"91",x"B2", -- 0x1488
    x"98",x"85",x"A6",x"18",x"60",x"A5",x"B9",x"30", -- 0x1490
    x"2C",x"A4",x"B7",x"F0",x"28",x"A5",x"BA",x"20", -- 0x1498
    x"17",x"EE",x"A5",x"B9",x"09",x"F0",x"20",x"C0", -- 0x14A0
    x"EE",x"A5",x"90",x"10",x"05",x"68",x"68",x"4C", -- 0x14A8
    x"8A",x"F7",x"A5",x"B7",x"F0",x"0C",x"A0",x"00", -- 0x14B0
    x"B1",x"BB",x"20",x"E4",x"EE",x"C8",x"C4",x"B7", -- 0x14B8
    x"D0",x"F6",x"20",x"04",x"EF",x"18",x"60",x"A9", -- 0x14C0
    x"06",x"8D",x"12",x"91",x"8D",x"10",x"91",x"A9", -- 0x14C8
    x"EE",x"8D",x"1C",x"91",x"A0",x"00",x"8C",x"97", -- 0x14D0
    x"02",x"C4",x"B7",x"F0",x"0A",x"B1",x"BB",x"99", -- 0x14D8
    x"93",x"02",x"C8",x"C0",x"04",x"D0",x"F2",x"20", -- 0x14E0
    x"27",x"F0",x"8E",x"98",x"02",x"AD",x"93",x"02", -- 0x14E8
    x"29",x"0F",x"D0",x"00",x"0A",x"AA",x"BD",x"5A", -- 0x14F0
    x"FF",x"0A",x"A8",x"BD",x"5B",x"FF",x"2A",x"48", -- 0x14F8
    x"98",x"69",x"C8",x"8D",x"99",x"02",x"68",x"69", -- 0x1500
    x"00",x"8D",x"9A",x"02",x"AD",x"94",x"02",x"4A", -- 0x1508
    x"90",x"09",x"AD",x"20",x"91",x"0A",x"B0",x"03", -- 0x1510
    x"4C",x"16",x"F0",x"AD",x"9B",x"02",x"8D",x"9C", -- 0x1518
    x"02",x"AD",x"9E",x"02",x"8D",x"9D",x"02",x"20", -- 0x1520
    x"75",x"FE",x"A5",x"F8",x"D0",x"05",x"88",x"84", -- 0x1528
    x"F8",x"86",x"F7",x"A5",x"FA",x"D0",x"05",x"88", -- 0x1530
    x"84",x"FA",x"86",x"F9",x"38",x"A9",x"F0",x"4C", -- 0x1538
    x"7B",x"FE",x"86",x"C3",x"84",x"C4",x"6C",x"30", -- 0x1540
    x"03",x"85",x"93",x"A9",x"00",x"85",x"90",x"A5", -- 0x1548
    x"BA",x"D0",x"03",x"4C",x"96",x"F7",x"C9",x"03", -- 0x1550
    x"F0",x"F9",x"90",x"6E",x"A4",x"B7",x"D0",x"03", -- 0x1558
    x"4C",x"93",x"F7",x"20",x"BC",x"E4",x"A9",x"60", -- 0x1560
    x"85",x"B9",x"20",x"95",x"F4",x"A5",x"BA",x"20", -- 0x1568
    x"14",x"EE",x"A5",x"B9",x"20",x"CE",x"EE",x"20", -- 0x1570
    x"19",x"EF",x"85",x"AE",x"A5",x"90",x"4A",x"4A", -- 0x1578
    x"B0",x"45",x"20",x"19",x"EF",x"85",x"AF",x"20", -- 0x1580
    x"C1",x"E4",x"A9",x"FD",x"25",x"90",x"85",x"90", -- 0x1588
    x"20",x"E1",x"FF",x"D0",x"03",x"4C",x"CB",x"F6", -- 0x1590
    x"20",x"19",x"EF",x"AA",x"A5",x"90",x"4A",x"4A", -- 0x1598
    x"B0",x"E8",x"8A",x"A4",x"93",x"F0",x"0C",x"A0", -- 0x15A0
    x"00",x"D1",x"AE",x"F0",x"08",x"A9",x"10",x"20", -- 0x15A8
    x"6A",x"FE",x"2C",x"91",x"AE",x"E6",x"AE",x"D0", -- 0x15B0
    x"02",x"E6",x"AF",x"24",x"90",x"50",x"CB",x"20", -- 0x15B8
    x"F6",x"EE",x"20",x"DA",x"F6",x"90",x"7A",x"4C", -- 0x15C0
    x"87",x"F7",x"C9",x"02",x"D0",x"03",x"4C",x"B9", -- 0x15C8
    x"F0",x"20",x"4D",x"F8",x"B0",x"03",x"4C",x"96", -- 0x15D0
    x"F7",x"20",x"94",x"F8",x"B0",x"68",x"20",x"47", -- 0x15D8
    x"F6",x"A5",x"B7",x"F0",x"09",x"20",x"67",x"F8", -- 0x15E0
    x"90",x"0B",x"F0",x"5A",x"B0",x"D9",x"20",x"AF", -- 0x15E8
    x"F7",x"F0",x"53",x"B0",x"D2",x"A5",x"90",x"29", -- 0x15F0
    x"10",x"38",x"D0",x"4A",x"E0",x"01",x"F0",x"11", -- 0x15F8
    x"E0",x"03",x"D0",x"DD",x"A0",x"01",x"B1",x"B2", -- 0x1600
    x"85",x"C3",x"C8",x"B1",x"B2",x"85",x"C4",x"B0", -- 0x1608
    x"04",x"A5",x"B9",x"D0",x"EF",x"A0",x"03",x"B1", -- 0x1610
    x"B2",x"A0",x"01",x"F1",x"B2",x"AA",x"A0",x"04", -- 0x1618
    x"B1",x"B2",x"A0",x"02",x"F1",x"B2",x"A8",x"18", -- 0x1620
    x"8A",x"65",x"C3",x"85",x"AE",x"98",x"65",x"C4", -- 0x1628
    x"85",x"AF",x"A5",x"C3",x"85",x"C1",x"A5",x"C4", -- 0x1630
    x"85",x"C2",x"20",x"6A",x"F6",x"20",x"C9",x"F8", -- 0x1638
    x"24",x"18",x"A6",x"AE",x"A4",x"AF",x"60",x"A5", -- 0x1640
    x"9D",x"10",x"1E",x"A0",x"0C",x"20",x"E6",x"F1", -- 0x1648
    x"A5",x"B7",x"F0",x"15",x"A0",x"17",x"20",x"E6", -- 0x1650
    x"F1",x"A4",x"B7",x"F0",x"0C",x"A0",x"00",x"B1", -- 0x1658
    x"BB",x"20",x"D2",x"FF",x"C8",x"C4",x"B7",x"D0", -- 0x1660
    x"F6",x"60",x"A0",x"49",x"A5",x"93",x"F0",x"02", -- 0x1668
    x"A0",x"59",x"4C",x"E2",x"F1",x"86",x"AE",x"84", -- 0x1670
    x"AF",x"AA",x"B5",x"00",x"85",x"C1",x"B5",x"01", -- 0x1678
    x"85",x"C2",x"6C",x"32",x"03",x"A5",x"BA",x"D0", -- 0x1680
    x"03",x"4C",x"96",x"F7",x"C9",x"03",x"F0",x"F9", -- 0x1688
    x"90",x"5F",x"A9",x"61",x"85",x"B9",x"A4",x"B7", -- 0x1690
    x"D0",x"03",x"4C",x"93",x"F7",x"20",x"95",x"F4", -- 0x1698
    x"20",x"28",x"F7",x"A5",x"BA",x"20",x"17",x"EE", -- 0x16A0
    x"A5",x"B9",x"20",x"C0",x"EE",x"A0",x"00",x"20", -- 0x16A8
    x"D2",x"FB",x"A5",x"AC",x"20",x"E4",x"EE",x"A5", -- 0x16B0
    x"AD",x"20",x"E4",x"EE",x"20",x"11",x"FD",x"B0", -- 0x16B8
    x"16",x"B1",x"AC",x"20",x"E4",x"EE",x"20",x"E1", -- 0x16C0
    x"FF",x"D0",x"07",x"20",x"DA",x"F6",x"A9",x"00", -- 0x16C8
    x"38",x"60",x"20",x"1B",x"FD",x"D0",x"E5",x"20", -- 0x16D0
    x"04",x"EF",x"24",x"B9",x"30",x"11",x"A5",x"BA", -- 0x16D8
    x"20",x"17",x"EE",x"A5",x"B9",x"29",x"EF",x"09", -- 0x16E0
    x"E0",x"20",x"C0",x"EE",x"20",x"04",x"EF",x"18", -- 0x16E8
    x"60",x"C9",x"02",x"D0",x"03",x"4C",x"B9",x"F0", -- 0x16F0
    x"20",x"4D",x"F8",x"90",x"8C",x"20",x"B7",x"F8", -- 0x16F8
    x"B0",x"25",x"20",x"28",x"F7",x"A2",x"03",x"A5", -- 0x1700
    x"B9",x"29",x"01",x"D0",x"02",x"A2",x"01",x"8A", -- 0x1708
    x"20",x"E7",x"F7",x"B0",x"12",x"20",x"E6",x"F8", -- 0x1710
    x"B0",x"0D",x"A5",x"B9",x"29",x"02",x"F0",x"06", -- 0x1718
    x"A9",x"05",x"20",x"E7",x"F7",x"24",x"18",x"60", -- 0x1720
    x"A5",x"9D",x"10",x"FB",x"A0",x"51",x"20",x"E6", -- 0x1728
    x"F1",x"4C",x"59",x"F6",x"A2",x"00",x"E6",x"A2", -- 0x1730
    x"D0",x"06",x"E6",x"A1",x"D0",x"02",x"E6",x"A0", -- 0x1738
    x"38",x"A5",x"A2",x"E9",x"01",x"A5",x"A1",x"E9", -- 0x1740
    x"1A",x"A5",x"A0",x"E9",x"4F",x"90",x"06",x"86", -- 0x1748
    x"A0",x"86",x"A1",x"86",x"A2",x"AD",x"2F",x"91", -- 0x1750
    x"CD",x"2F",x"91",x"D0",x"F8",x"85",x"91",x"60", -- 0x1758
    x"78",x"A5",x"A2",x"A6",x"A1",x"A4",x"A0",x"78", -- 0x1760
    x"85",x"A2",x"86",x"A1",x"84",x"A0",x"58",x"60", -- 0x1768
    x"A5",x"91",x"C9",x"FE",x"D0",x"07",x"08",x"20", -- 0x1770
    x"CC",x"FF",x"85",x"C6",x"28",x"60",x"A9",x"01", -- 0x1778
    x"2C",x"A9",x"02",x"2C",x"A9",x"03",x"2C",x"A9", -- 0x1780
    x"04",x"2C",x"A9",x"05",x"2C",x"A9",x"06",x"2C", -- 0x1788
    x"A9",x"07",x"2C",x"A9",x"08",x"2C",x"A9",x"09", -- 0x1790
    x"48",x"20",x"CC",x"FF",x"A0",x"00",x"24",x"9D", -- 0x1798
    x"50",x"0A",x"20",x"E6",x"F1",x"68",x"48",x"09", -- 0x17A0
    x"30",x"20",x"D2",x"FF",x"68",x"38",x"60",x"A5", -- 0x17A8
    x"93",x"48",x"20",x"C0",x"F8",x"68",x"85",x"93", -- 0x17B0
    x"B0",x"2C",x"A0",x"00",x"B1",x"B2",x"C9",x"05", -- 0x17B8
    x"F0",x"24",x"C9",x"01",x"F0",x"08",x"C9",x"03", -- 0x17C0
    x"F0",x"04",x"C9",x"04",x"D0",x"E1",x"AA",x"24", -- 0x17C8
    x"9D",x"10",x"11",x"A0",x"63",x"20",x"E6",x"F1", -- 0x17D0
    x"A0",x"05",x"B1",x"B2",x"20",x"D2",x"FF",x"C8", -- 0x17D8
    x"C0",x"15",x"D0",x"F6",x"18",x"88",x"60",x"85", -- 0x17E0
    x"9E",x"20",x"4D",x"F8",x"90",x"5E",x"A5",x"C2", -- 0x17E8
    x"48",x"A5",x"C1",x"48",x"A5",x"AF",x"48",x"A5", -- 0x17F0
    x"AE",x"48",x"A0",x"BF",x"A9",x"20",x"91",x"B2", -- 0x17F8
    x"88",x"D0",x"FB",x"A5",x"9E",x"91",x"B2",x"C8", -- 0x1800
    x"A5",x"C1",x"91",x"B2",x"C8",x"A5",x"C2",x"91", -- 0x1808
    x"B2",x"C8",x"A5",x"AE",x"91",x"B2",x"C8",x"A5", -- 0x1810
    x"AF",x"91",x"B2",x"C8",x"84",x"9F",x"A0",x"00", -- 0x1818
    x"84",x"9E",x"A4",x"9E",x"C4",x"B7",x"F0",x"0C", -- 0x1820
    x"B1",x"BB",x"A4",x"9F",x"91",x"B2",x"E6",x"9E", -- 0x1828
    x"E6",x"9F",x"D0",x"EE",x"20",x"54",x"F8",x"A9", -- 0x1830
    x"69",x"85",x"AB",x"20",x"EA",x"F8",x"A8",x"68", -- 0x1838
    x"85",x"AE",x"68",x"85",x"AF",x"68",x"85",x"C1", -- 0x1840
    x"68",x"85",x"C2",x"98",x"60",x"A6",x"B2",x"A4", -- 0x1848
    x"B3",x"C0",x"02",x"60",x"20",x"4D",x"F8",x"8A", -- 0x1850
    x"85",x"C1",x"18",x"69",x"C0",x"85",x"AE",x"98", -- 0x1858
    x"85",x"C2",x"69",x"00",x"85",x"AF",x"60",x"20", -- 0x1860
    x"AF",x"F7",x"B0",x"1D",x"A0",x"05",x"84",x"9F", -- 0x1868
    x"A0",x"00",x"84",x"9E",x"C4",x"B7",x"F0",x"10", -- 0x1870
    x"B1",x"BB",x"A4",x"9F",x"D1",x"B2",x"D0",x"E7", -- 0x1878
    x"E6",x"9E",x"E6",x"9F",x"A4",x"9E",x"D0",x"EC", -- 0x1880
    x"18",x"60",x"20",x"4D",x"F8",x"E6",x"A6",x"A4", -- 0x1888
    x"A6",x"C0",x"C0",x"60",x"20",x"AB",x"F8",x"F0", -- 0x1890
    x"1C",x"A0",x"1B",x"20",x"E6",x"F1",x"20",x"4B", -- 0x1898
    x"F9",x"20",x"AB",x"F8",x"D0",x"F8",x"A0",x"6A", -- 0x18A0
    x"4C",x"E6",x"F1",x"A9",x"40",x"2C",x"1F",x"91", -- 0x18A8
    x"D0",x"03",x"2C",x"1F",x"91",x"18",x"60",x"20", -- 0x18B0
    x"AB",x"F8",x"F0",x"F9",x"A0",x"2E",x"D0",x"DB", -- 0x18B8
    x"A9",x"00",x"85",x"90",x"85",x"93",x"20",x"54", -- 0x18C0
    x"F8",x"20",x"94",x"F8",x"B0",x"1F",x"78",x"A9", -- 0x18C8
    x"00",x"85",x"AA",x"85",x"B4",x"85",x"B0",x"85", -- 0x18D0
    x"9E",x"85",x"9F",x"85",x"9C",x"A9",x"82",x"A2", -- 0x18D8
    x"0E",x"D0",x"11",x"20",x"54",x"F8",x"A9",x"14", -- 0x18E0
    x"85",x"AB",x"20",x"B7",x"F8",x"B0",x"68",x"78", -- 0x18E8
    x"A9",x"A0",x"A2",x"08",x"A0",x"7F",x"8C",x"2E", -- 0x18F0
    x"91",x"8D",x"2E",x"91",x"20",x"60",x"F1",x"AD", -- 0x18F8
    x"14",x"03",x"8D",x"9F",x"02",x"AD",x"15",x"03", -- 0x1900
    x"8D",x"A0",x"02",x"20",x"FB",x"FC",x"A9",x"02", -- 0x1908
    x"85",x"BE",x"20",x"DB",x"FB",x"AD",x"1C",x"91", -- 0x1910
    x"29",x"FD",x"09",x"0C",x"8D",x"1C",x"91",x"85", -- 0x1918
    x"C0",x"A2",x"FF",x"A0",x"FF",x"88",x"D0",x"FD", -- 0x1920
    x"CA",x"D0",x"F8",x"8D",x"29",x"91",x"58",x"AD", -- 0x1928
    x"A0",x"02",x"CD",x"15",x"03",x"18",x"F0",x"1F", -- 0x1930
    x"20",x"4B",x"F9",x"AD",x"2D",x"91",x"29",x"40", -- 0x1938
    x"F0",x"ED",x"AD",x"14",x"91",x"20",x"34",x"F7", -- 0x1940
    x"4C",x"2F",x"F9",x"20",x"E1",x"FF",x"18",x"D0", -- 0x1948
    x"0B",x"20",x"CF",x"FC",x"38",x"68",x"68",x"A9", -- 0x1950
    x"00",x"8D",x"A0",x"02",x"60",x"86",x"B1",x"A5", -- 0x1958
    x"B0",x"0A",x"0A",x"18",x"65",x"B0",x"18",x"65", -- 0x1960
    x"B1",x"85",x"B1",x"A9",x"00",x"24",x"B0",x"30", -- 0x1968
    x"01",x"2A",x"06",x"B1",x"2A",x"06",x"B1",x"2A", -- 0x1970
    x"AA",x"AD",x"28",x"91",x"C9",x"15",x"90",x"F9", -- 0x1978
    x"65",x"B1",x"8D",x"24",x"91",x"8A",x"6D",x"29", -- 0x1980
    x"91",x"8D",x"25",x"91",x"58",x"60",x"AE",x"29", -- 0x1988
    x"91",x"A0",x"FF",x"98",x"ED",x"28",x"91",x"EC", -- 0x1990
    x"29",x"91",x"D0",x"F2",x"86",x"B1",x"AA",x"8C", -- 0x1998
    x"28",x"91",x"8C",x"29",x"91",x"98",x"E5",x"B1", -- 0x19A0
    x"86",x"B1",x"4A",x"66",x"B1",x"4A",x"66",x"B1", -- 0x19A8
    x"A5",x"B0",x"18",x"69",x"3C",x"2C",x"21",x"91", -- 0x19B0
    x"C5",x"B1",x"B0",x"4A",x"A6",x"9C",x"F0",x"03", -- 0x19B8
    x"4C",x"AD",x"FA",x"A6",x"A3",x"30",x"1B",x"A2", -- 0x19C0
    x"00",x"69",x"30",x"65",x"B0",x"C5",x"B1",x"B0", -- 0x19C8
    x"1C",x"E8",x"69",x"26",x"65",x"B0",x"C5",x"B1", -- 0x19D0
    x"B0",x"17",x"69",x"2C",x"65",x"B0",x"C5",x"B1", -- 0x19D8
    x"90",x"03",x"4C",x"60",x"FA",x"A5",x"B4",x"F0", -- 0x19E0
    x"1D",x"85",x"A8",x"D0",x"19",x"E6",x"A9",x"B0", -- 0x19E8
    x"02",x"C6",x"A9",x"38",x"E9",x"13",x"E5",x"B1", -- 0x19F0
    x"65",x"92",x"85",x"92",x"A5",x"A4",x"49",x"01", -- 0x19F8
    x"85",x"A4",x"F0",x"21",x"86",x"D7",x"A5",x"B4", -- 0x1A00
    x"F0",x"18",x"2C",x"2D",x"91",x"50",x"13",x"A9", -- 0x1A08
    x"00",x"85",x"A4",x"A5",x"A3",x"10",x"30",x"30", -- 0x1A10
    x"C9",x"A2",x"A6",x"20",x"5D",x"F9",x"A5",x"9B", -- 0x1A18
    x"D0",x"C3",x"4C",x"56",x"FF",x"A5",x"92",x"F0", -- 0x1A20
    x"07",x"30",x"03",x"C6",x"B0",x"2C",x"E6",x"B0", -- 0x1A28
    x"A9",x"00",x"85",x"92",x"E4",x"D7",x"D0",x"0F", -- 0x1A30
    x"8A",x"D0",x"AA",x"A5",x"A9",x"30",x"C7",x"C9", -- 0x1A38
    x"10",x"90",x"C3",x"85",x"96",x"B0",x"BF",x"8A", -- 0x1A40
    x"45",x"9B",x"85",x"9B",x"A5",x"B4",x"F0",x"D2", -- 0x1A48
    x"C6",x"A3",x"30",x"C5",x"46",x"D7",x"66",x"BF", -- 0x1A50
    x"A2",x"DA",x"20",x"5D",x"F9",x"4C",x"56",x"FF", -- 0x1A58
    x"A5",x"96",x"F0",x"04",x"A5",x"B4",x"F0",x"04", -- 0x1A60
    x"A5",x"A3",x"10",x"85",x"46",x"B1",x"A9",x"93", -- 0x1A68
    x"38",x"E5",x"B1",x"65",x"B0",x"0A",x"AA",x"20", -- 0x1A70
    x"5D",x"F9",x"E6",x"9C",x"A5",x"B4",x"D0",x"11", -- 0x1A78
    x"A5",x"96",x"F0",x"26",x"85",x"A8",x"A9",x"00", -- 0x1A80
    x"85",x"96",x"A9",x"C0",x"8D",x"2E",x"91",x"85", -- 0x1A88
    x"B4",x"A5",x"96",x"85",x"B5",x"F0",x"09",x"A9", -- 0x1A90
    x"00",x"85",x"B4",x"A9",x"40",x"8D",x"2E",x"91", -- 0x1A98
    x"A5",x"BF",x"85",x"BD",x"A5",x"A8",x"05",x"A9", -- 0x1AA0
    x"85",x"B6",x"4C",x"56",x"FF",x"20",x"DB",x"FB", -- 0x1AA8
    x"85",x"9C",x"A2",x"DA",x"20",x"5D",x"F9",x"A5", -- 0x1AB0
    x"BE",x"F0",x"02",x"85",x"A7",x"A9",x"0F",x"24", -- 0x1AB8
    x"AA",x"10",x"17",x"A5",x"B5",x"D0",x"0C",x"A6", -- 0x1AC0
    x"BE",x"CA",x"D0",x"0B",x"A9",x"08",x"20",x"6A", -- 0x1AC8
    x"FE",x"D0",x"04",x"A9",x"00",x"85",x"AA",x"4C", -- 0x1AD0
    x"56",x"FF",x"70",x"31",x"D0",x"18",x"A5",x"B5", -- 0x1AD8
    x"D0",x"F5",x"A5",x"B6",x"D0",x"F1",x"A5",x"A7", -- 0x1AE0
    x"4A",x"A5",x"BD",x"30",x"03",x"90",x"18",x"18", -- 0x1AE8
    x"B0",x"15",x"29",x"0F",x"85",x"AA",x"C6",x"AA", -- 0x1AF0
    x"D0",x"DD",x"A9",x"40",x"85",x"AA",x"20",x"D2", -- 0x1AF8
    x"FB",x"A9",x"00",x"85",x"AB",x"F0",x"D0",x"A9", -- 0x1B00
    x"80",x"85",x"AA",x"D0",x"CA",x"A5",x"B5",x"F0", -- 0x1B08
    x"0A",x"A9",x"04",x"20",x"6A",x"FE",x"A9",x"00", -- 0x1B10
    x"4C",x"97",x"FB",x"20",x"11",x"FD",x"90",x"03", -- 0x1B18
    x"4C",x"95",x"FB",x"A6",x"A7",x"CA",x"F0",x"2D", -- 0x1B20
    x"A5",x"93",x"F0",x"0C",x"A0",x"00",x"A5",x"BD", -- 0x1B28
    x"D1",x"AC",x"F0",x"04",x"A9",x"01",x"85",x"B6", -- 0x1B30
    x"A5",x"B6",x"F0",x"4B",x"A2",x"3D",x"E4",x"9E", -- 0x1B38
    x"90",x"3E",x"A6",x"9E",x"A5",x"AD",x"9D",x"01", -- 0x1B40
    x"01",x"A5",x"AC",x"9D",x"00",x"01",x"E8",x"E8", -- 0x1B48
    x"86",x"9E",x"4C",x"87",x"FB",x"A6",x"9F",x"E4", -- 0x1B50
    x"9E",x"F0",x"35",x"A5",x"AC",x"DD",x"00",x"01", -- 0x1B58
    x"D0",x"2E",x"A5",x"AD",x"DD",x"01",x"01",x"D0", -- 0x1B60
    x"27",x"E6",x"9F",x"E6",x"9F",x"A5",x"93",x"F0", -- 0x1B68
    x"0B",x"A5",x"BD",x"A0",x"00",x"D1",x"AC",x"F0", -- 0x1B70
    x"17",x"C8",x"84",x"B6",x"A5",x"B6",x"F0",x"07", -- 0x1B78
    x"A9",x"10",x"20",x"6A",x"FE",x"D0",x"09",x"A5", -- 0x1B80
    x"93",x"D0",x"05",x"A8",x"A5",x"BD",x"91",x"AC", -- 0x1B88
    x"20",x"1B",x"FD",x"D0",x"3A",x"A9",x"80",x"85", -- 0x1B90
    x"AA",x"A6",x"BE",x"CA",x"30",x"02",x"86",x"BE", -- 0x1B98
    x"C6",x"A7",x"F0",x"08",x"A5",x"9E",x"D0",x"27", -- 0x1BA0
    x"85",x"BE",x"F0",x"23",x"20",x"CF",x"FC",x"20", -- 0x1BA8
    x"D2",x"FB",x"A0",x"00",x"84",x"AB",x"B1",x"AC", -- 0x1BB0
    x"45",x"AB",x"85",x"AB",x"20",x"1B",x"FD",x"20", -- 0x1BB8
    x"11",x"FD",x"90",x"F2",x"A5",x"AB",x"45",x"BD", -- 0x1BC0
    x"F0",x"05",x"A9",x"20",x"20",x"6A",x"FE",x"4C", -- 0x1BC8
    x"56",x"FF",x"A5",x"C2",x"85",x"AD",x"A5",x"C1", -- 0x1BD0
    x"85",x"AC",x"60",x"A9",x"08",x"85",x"A3",x"A9", -- 0x1BD8
    x"00",x"85",x"A4",x"85",x"A8",x"85",x"9B",x"85", -- 0x1BE0
    x"A9",x"60",x"A5",x"BD",x"4A",x"A9",x"60",x"90", -- 0x1BE8
    x"02",x"A9",x"B0",x"A2",x"00",x"8D",x"28",x"91", -- 0x1BF0
    x"8E",x"29",x"91",x"AD",x"20",x"91",x"49",x"08", -- 0x1BF8
    x"8D",x"20",x"91",x"29",x"08",x"60",x"38",x"66", -- 0x1C00
    x"AD",x"30",x"3C",x"A5",x"A8",x"D0",x"12",x"A9", -- 0x1C08
    x"10",x"A2",x"01",x"20",x"F5",x"FB",x"D0",x"2F", -- 0x1C10
    x"E6",x"A8",x"A5",x"AD",x"10",x"29",x"4C",x"95", -- 0x1C18
    x"FC",x"A5",x"A9",x"D0",x"09",x"20",x"F1",x"FB", -- 0x1C20
    x"D0",x"1D",x"E6",x"A9",x"D0",x"19",x"20",x"EA", -- 0x1C28
    x"FB",x"D0",x"14",x"A5",x"A4",x"49",x"01",x"85", -- 0x1C30
    x"A4",x"F0",x"0F",x"A5",x"BD",x"49",x"01",x"85", -- 0x1C38
    x"BD",x"29",x"01",x"45",x"9B",x"85",x"9B",x"4C", -- 0x1C40
    x"56",x"FF",x"46",x"BD",x"C6",x"A3",x"A5",x"A3", -- 0x1C48
    x"F0",x"3A",x"10",x"F3",x"20",x"DB",x"FB",x"58", -- 0x1C50
    x"A5",x"A5",x"F0",x"12",x"A2",x"00",x"86",x"D7", -- 0x1C58
    x"C6",x"A5",x"A6",x"BE",x"E0",x"02",x"D0",x"02", -- 0x1C60
    x"09",x"80",x"85",x"BD",x"D0",x"D9",x"20",x"11", -- 0x1C68
    x"FD",x"90",x"0A",x"D0",x"91",x"E6",x"AD",x"A5", -- 0x1C70
    x"D7",x"85",x"BD",x"B0",x"CA",x"A0",x"00",x"B1", -- 0x1C78
    x"AC",x"85",x"BD",x"45",x"D7",x"85",x"D7",x"20", -- 0x1C80
    x"1B",x"FD",x"D0",x"BB",x"A5",x"9B",x"49",x"01", -- 0x1C88
    x"85",x"BD",x"4C",x"56",x"FF",x"C6",x"BE",x"D0", -- 0x1C90
    x"03",x"20",x"08",x"FD",x"A9",x"50",x"85",x"A7", -- 0x1C98
    x"A2",x"08",x"78",x"20",x"FB",x"FC",x"D0",x"EA", -- 0x1CA0
    x"A9",x"78",x"20",x"F3",x"FB",x"D0",x"E3",x"C6", -- 0x1CA8
    x"A7",x"D0",x"DF",x"20",x"DB",x"FB",x"C6",x"AB", -- 0x1CB0
    x"10",x"D8",x"A2",x"0A",x"20",x"FB",x"FC",x"58", -- 0x1CB8
    x"E6",x"AB",x"A5",x"BE",x"F0",x"30",x"20",x"D2", -- 0x1CC0
    x"FB",x"A2",x"09",x"86",x"A5",x"D0",x"85",x"08", -- 0x1CC8
    x"78",x"20",x"08",x"FD",x"A9",x"7F",x"8D",x"2E", -- 0x1CD0
    x"91",x"A9",x"F7",x"8D",x"20",x"91",x"A9",x"40", -- 0x1CD8
    x"8D",x"2B",x"91",x"20",x"39",x"FE",x"AD",x"A0", -- 0x1CE0
    x"02",x"F0",x"09",x"8D",x"15",x"03",x"AD",x"9F", -- 0x1CE8
    x"02",x"8D",x"14",x"03",x"28",x"60",x"20",x"CF", -- 0x1CF0
    x"FC",x"F0",x"97",x"BD",x"E9",x"FD",x"8D",x"14", -- 0x1CF8
    x"03",x"BD",x"EA",x"FD",x"8D",x"15",x"03",x"60", -- 0x1D00
    x"AD",x"1C",x"91",x"09",x"0E",x"8D",x"1C",x"91", -- 0x1D08
    x"60",x"38",x"A5",x"AC",x"E5",x"AE",x"A5",x"AD", -- 0x1D10
    x"E5",x"AF",x"60",x"E6",x"AC",x"D0",x"02",x"E6", -- 0x1D18
    x"AD",x"60",x"A2",x"FF",x"78",x"9A",x"D8",x"20", -- 0x1D20
    x"3F",x"FD",x"D0",x"03",x"6C",x"00",x"A0",x"20", -- 0x1D28
    x"8D",x"FD",x"20",x"52",x"FD",x"20",x"F9",x"FD", -- 0x1D30
    x"20",x"18",x"E5",x"58",x"6C",x"00",x"C0",x"A2", -- 0x1D38
    x"05",x"BD",x"4C",x"FD",x"DD",x"03",x"A0",x"D0", -- 0x1D40
    x"03",x"CA",x"D0",x"F5",x"60",x"41",x"30",x"C3", -- 0x1D48
    x"C2",x"CD",x"A2",x"6D",x"A0",x"FD",x"18",x"86", -- 0x1D50
    x"C3",x"84",x"C4",x"A0",x"1F",x"B9",x"14",x"03", -- 0x1D58
    x"B0",x"02",x"B1",x"C3",x"91",x"C3",x"99",x"14", -- 0x1D60
    x"03",x"88",x"10",x"F1",x"60",x"BF",x"EA",x"D2", -- 0x1D68
    x"FE",x"AD",x"FE",x"0A",x"F4",x"4A",x"F3",x"C7", -- 0x1D70
    x"F2",x"09",x"F3",x"F3",x"F3",x"0E",x"F2",x"7A", -- 0x1D78
    x"F2",x"70",x"F7",x"F5",x"F1",x"EF",x"F3",x"D2", -- 0x1D80
    x"FE",x"49",x"F5",x"85",x"F6",x"A9",x"00",x"AA", -- 0x1D88
    x"95",x"00",x"9D",x"00",x"02",x"9D",x"00",x"03", -- 0x1D90
    x"E8",x"D0",x"F5",x"A2",x"3C",x"A0",x"03",x"86", -- 0x1D98
    x"B2",x"84",x"B3",x"85",x"C1",x"85",x"97",x"8D", -- 0x1DA0
    x"81",x"02",x"A8",x"A9",x"04",x"85",x"C2",x"E6", -- 0x1DA8
    x"C1",x"D0",x"02",x"E6",x"C2",x"20",x"91",x"FE", -- 0x1DB0
    x"A5",x"97",x"F0",x"22",x"B0",x"F1",x"A4",x"C2", -- 0x1DB8
    x"A6",x"C1",x"C0",x"20",x"90",x"25",x"C0",x"21", -- 0x1DC0
    x"B0",x"08",x"A0",x"1E",x"8C",x"88",x"02",x"4C", -- 0x1DC8
    x"7B",x"FE",x"A9",x"12",x"8D",x"82",x"02",x"A9", -- 0x1DD0
    x"10",x"8D",x"88",x"02",x"D0",x"F1",x"90",x"CF", -- 0x1DD8
    x"A5",x"C2",x"8D",x"82",x"02",x"85",x"97",x"C9", -- 0x1DE0
    x"11",x"90",x"C4",x"20",x"C3",x"E5",x"4C",x"EB", -- 0x1DE8
    x"FD",x"A8",x"FC",x"0B",x"FC",x"BF",x"EA",x"8E", -- 0x1DF0
    x"F9",x"A9",x"7F",x"8D",x"1E",x"91",x"8D",x"2E", -- 0x1DF8
    x"91",x"A9",x"40",x"8D",x"2B",x"91",x"A9",x"40", -- 0x1E00
    x"8D",x"1B",x"91",x"A9",x"FE",x"8D",x"1C",x"91", -- 0x1E08
    x"A9",x"DE",x"8D",x"2C",x"91",x"A2",x"00",x"8E", -- 0x1E10
    x"12",x"91",x"A2",x"FF",x"8E",x"22",x"91",x"A2", -- 0x1E18
    x"00",x"8E",x"23",x"91",x"A2",x"80",x"8E",x"13", -- 0x1E20
    x"91",x"A2",x"00",x"8E",x"1F",x"91",x"20",x"84", -- 0x1E28
    x"EF",x"A9",x"82",x"8D",x"1E",x"91",x"20",x"8D", -- 0x1E30
    x"EF",x"A9",x"C0",x"8D",x"2E",x"91",x"A9",x"26", -- 0x1E38
    x"8D",x"24",x"91",x"A9",x"48",x"8D",x"25",x"91", -- 0x1E40
    x"60",x"85",x"B7",x"86",x"BB",x"84",x"BC",x"60", -- 0x1E48
    x"85",x"B8",x"86",x"BA",x"84",x"B9",x"60",x"A5", -- 0x1E50
    x"BA",x"C9",x"02",x"D0",x"0B",x"AD",x"97",x"02", -- 0x1E58
    x"A9",x"00",x"8D",x"97",x"02",x"60",x"85",x"9D", -- 0x1E60
    x"A5",x"90",x"05",x"90",x"85",x"90",x"60",x"8D", -- 0x1E68
    x"85",x"02",x"60",x"90",x"06",x"AE",x"83",x"02", -- 0x1E70
    x"AC",x"84",x"02",x"8E",x"83",x"02",x"8C",x"84", -- 0x1E78
    x"02",x"60",x"90",x"06",x"AE",x"81",x"02",x"AC", -- 0x1E80
    x"82",x"02",x"8E",x"81",x"02",x"8C",x"82",x"02", -- 0x1E88
    x"60",x"B1",x"C1",x"AA",x"A9",x"55",x"91",x"C1", -- 0x1E90
    x"D1",x"C1",x"D0",x"08",x"6A",x"91",x"C1",x"D1", -- 0x1E98
    x"C1",x"D0",x"01",x"A9",x"18",x"8A",x"91",x"C1", -- 0x1EA0
    x"60",x"78",x"6C",x"18",x"03",x"48",x"8A",x"48", -- 0x1EA8
    x"98",x"48",x"AD",x"1D",x"91",x"10",x"48",x"2D", -- 0x1EB0
    x"1E",x"91",x"AA",x"29",x"02",x"F0",x"1F",x"20", -- 0x1EB8
    x"3F",x"FD",x"D0",x"03",x"6C",x"02",x"A0",x"2C", -- 0x1EC0
    x"11",x"91",x"20",x"34",x"F7",x"20",x"E1",x"FF", -- 0x1EC8
    x"D0",x"2D",x"20",x"52",x"FD",x"20",x"F9",x"FD", -- 0x1ED0
    x"20",x"18",x"E5",x"6C",x"02",x"C0",x"AD",x"1E", -- 0x1ED8
    x"91",x"09",x"80",x"48",x"A9",x"7F",x"8D",x"1E", -- 0x1EE0
    x"91",x"8A",x"29",x"40",x"F0",x"14",x"A9",x"CE", -- 0x1EE8
    x"05",x"B5",x"8D",x"1C",x"91",x"AD",x"14",x"91", -- 0x1EF0
    x"68",x"8D",x"1E",x"91",x"20",x"A3",x"EF",x"4C", -- 0x1EF8
    x"56",x"FF",x"8A",x"29",x"20",x"F0",x"25",x"AD", -- 0x1F00
    x"10",x"91",x"29",x"01",x"85",x"A7",x"AD",x"18", -- 0x1F08
    x"91",x"E9",x"16",x"6D",x"99",x"02",x"8D",x"18", -- 0x1F10
    x"91",x"AD",x"19",x"91",x"6D",x"9A",x"02",x"8D", -- 0x1F18
    x"19",x"91",x"68",x"8D",x"1E",x"91",x"20",x"36", -- 0x1F20
    x"F0",x"4C",x"56",x"FF",x"8A",x"29",x"10",x"F0", -- 0x1F28
    x"25",x"AD",x"93",x"02",x"29",x"0F",x"D0",x"00", -- 0x1F30
    x"0A",x"AA",x"BD",x"5A",x"FF",x"8D",x"18",x"91", -- 0x1F38
    x"BD",x"5B",x"FF",x"8D",x"19",x"91",x"AD",x"10", -- 0x1F40
    x"91",x"68",x"09",x"20",x"29",x"EF",x"8D",x"1E", -- 0x1F48
    x"91",x"AE",x"98",x"02",x"86",x"A8",x"68",x"A8", -- 0x1F50
    x"68",x"AA",x"68",x"40",x"E6",x"2A",x"78",x"1C", -- 0x1F58
    x"49",x"13",x"B1",x"0F",x"0A",x"0E",x"D3",x"06", -- 0x1F60
    x"38",x"03",x"6A",x"01",x"D0",x"00",x"83",x"00", -- 0x1F68
    x"36",x"00",x"48",x"8A",x"48",x"98",x"48",x"BA", -- 0x1F70
    x"BD",x"04",x"01",x"29",x"10",x"F0",x"03",x"6C", -- 0x1F78
    x"16",x"03",x"6C",x"14",x"03",x"FF",x"FF",x"FF", -- 0x1F80
    x"FF",x"FF",x"4C",x"52",x"FD",x"4C",x"57",x"FD", -- 0x1F88
    x"4C",x"66",x"FE",x"4C",x"C0",x"EE",x"4C",x"CE", -- 0x1F90
    x"EE",x"4C",x"73",x"FE",x"4C",x"82",x"FE",x"4C", -- 0x1F98
    x"1E",x"EB",x"4C",x"6F",x"FE",x"4C",x"19",x"EF", -- 0x1FA0
    x"4C",x"E4",x"EE",x"4C",x"F6",x"EE",x"4C",x"04", -- 0x1FA8
    x"EF",x"4C",x"17",x"EE",x"4C",x"14",x"EE",x"4C", -- 0x1FB0
    x"57",x"FE",x"4C",x"50",x"FE",x"4C",x"49",x"FE", -- 0x1FB8
    x"6C",x"1A",x"03",x"6C",x"1C",x"03",x"6C",x"1E", -- 0x1FC0
    x"03",x"6C",x"20",x"03",x"6C",x"22",x"03",x"6C", -- 0x1FC8
    x"24",x"03",x"6C",x"26",x"03",x"4C",x"42",x"F5", -- 0x1FD0
    x"4C",x"75",x"F6",x"4C",x"67",x"F7",x"4C",x"60", -- 0x1FD8
    x"F7",x"6C",x"28",x"03",x"6C",x"2A",x"03",x"6C", -- 0x1FE0
    x"2C",x"03",x"4C",x"34",x"F7",x"4C",x"05",x"E5", -- 0x1FE8
    x"4C",x"0A",x"E5",x"4C",x"00",x"E5",x"FF",x"FF", -- 0x1FF0
    x"FF",x"FF",x"A9",x"FE",x"22",x"FD",x"72",x"FF"  -- 0x1FF8
  );

begin

  p_rom : process
  begin
    wait until rising_edge(CLK);
     DATA <= ROM(to_integer(unsigned(ADDR)));
  end process;
end RTL;
