-------------------------------------------------------------------------------
-- $Id: vp_keymap-c.vhd,v 1.1 2007/02/10 12:53:52 arnim Exp $
-------------------------------------------------------------------------------

configuration vp_keymap_rtl_c0 of vp_keymap is

  for rtl
  end for;

end vp_keymap_rtl_c0;
