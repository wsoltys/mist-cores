
configuration key_slice_key_rom_c0 of key_slice is

  for key_rom
  end for;

end key_slice_key_rom_c0;
