-------------------------------------------------------------------------------
--
-- FPGA Videopac
--
-- $Id: rom_t48-c.vhd,v 1.2 2007/02/05 21:55:18 arnim Exp $
--
-------------------------------------------------------------------------------

configuration rom_t48_rtl_c0 of rom_t48 is

  for rtl
  end for;

end rom_t48_rtl_c0;
