-------------------------------------------------------------------------------
--
-- FPGA Videopac
--
-- $Id: vp_glue-c.vhd,v 1.4 2007/02/05 21:55:18 arnim Exp $
--
-------------------------------------------------------------------------------

configuration vp_glue_rtl_c0 of vp_glue is

  for rtl
  end for;

end vp_glue_rtl_c0;
