-- generated with romgen by MikeJ
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity rom_t48 is
  port (
    CLK         : in    std_logic;
    A           : in    std_logic_vector(9 downto 0);
    D           : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of rom_t48 is


  type ROM_ARRAY is array(0 to 1023) of std_logic_vector(7 downto 0);
  constant ROM : ROM_ARRAY := (
    x"84",x"00",x"00",x"84",x"02",x"00",x"00",x"84", -- 0x0000
    x"04",x"C5",x"AD",x"09",x"AE",x"14",x"E7",x"B8", -- 0x0008
    x"A1",x"80",x"72",x"18",x"FE",x"39",x"FD",x"93", -- 0x0010
    x"84",x"06",x"A5",x"B5",x"B9",x"A2",x"B8",x"3D", -- 0x0018
    x"81",x"A0",x"18",x"10",x"F0",x"53",x"3F",x"D3", -- 0x0020
    x"3C",x"96",x"2F",x"F0",x"53",x"C0",x"A0",x"18", -- 0x0028
    x"F0",x"37",x"F2",x"3A",x"37",x"53",x"7F",x"A0", -- 0x0030
    x"14",x"89",x"B9",x"3F",x"F1",x"37",x"D2",x"14", -- 0x0038
    x"EB",x"14",x"84",x"0A",x"FC",x"E3",x"A9",x"1C", -- 0x0040
    x"FC",x"E3",x"AA",x"F9",x"F2",x"5C",x"D2",x"73", -- 0x0048
    x"B2",x"7D",x"92",x"84",x"B9",x"3F",x"F1",x"53", -- 0x0050
    x"BF",x"A1",x"04",x"14",x"53",x"7F",x"AB",x"B8", -- 0x0058
    x"AA",x"27",x"90",x"B8",x"A7",x"B9",x"03",x"FA", -- 0x0060
    x"E3",x"90",x"18",x"1A",x"E9",x"67",x"FA",x"E3", -- 0x0068
    x"AA",x"04",x"76",x"53",x"3F",x"AB",x"1C",x"B8", -- 0x0070
    x"AA",x"FA",x"90",x"04",x"14",x"53",x"1F",x"AB", -- 0x0078
    x"BA",x"00",x"04",x"77",x"FA",x"AC",x"84",x"0A", -- 0x0080
    x"00",x"B8",x"7F",x"B9",x"A0",x"81",x"53",x"D6", -- 0x0088
    x"91",x"89",x"7C",x"99",x"E7",x"80",x"96",x"A3", -- 0x0090
    x"89",x"BC",x"99",x"B7",x"B9",x"A0",x"81",x"43", -- 0x0098
    x"28",x"91",x"83",x"AA",x"C8",x"80",x"A9",x"C8", -- 0x00A0
    x"80",x"91",x"C8",x"19",x"EA",x"A8",x"04",x"95", -- 0x00A8
    x"15",x"C5",x"09",x"AE",x"89",x"BC",x"99",x"BB", -- 0x00B0
    x"B8",x"F0",x"BA",x"06",x"F8",x"3A",x"0A",x"92", -- 0x00B8
    x"DA",x"BA",x"30",x"A8",x"0A",x"D8",x"96",x"DF", -- 0x00C0
    x"EA",x"C4",x"F8",x"47",x"77",x"D3",x"07",x"53", -- 0x00C8
    x"3F",x"A9",x"FF",x"53",x"3F",x"D9",x"96",x"E5", -- 0x00D0
    x"04",x"DF",x"18",x"EA",x"BC",x"BF",x"FF",x"FF", -- 0x00D8
    x"43",x"C0",x"AF",x"64",x"78",x"64",x"76",x"89", -- 0x00E0
    x"BC",x"99",x"B7",x"83",x"89",x"BC",x"99",x"AF", -- 0x00E8
    x"83",x"89",x"BC",x"99",x"B7",x"23",x"20",x"A8", -- 0x00F0
    x"A9",x"27",x"A0",x"18",x"E9",x"FA",x"14",x"EC", -- 0x00F8
    x"B9",x"FF",x"91",x"E9",x"02",x"91",x"14",x"E7", -- 0x0100
    x"34",x"1C",x"B8",x"FF",x"B9",x"80",x"27",x"90", -- 0x0108
    x"C8",x"E9",x"0F",x"23",x"F8",x"90",x"E8",x"15", -- 0x0110
    x"90",x"34",x"27",x"83",x"15",x"C5",x"B8",x"A0", -- 0x0118
    x"80",x"53",x"D6",x"90",x"D5",x"05",x"83",x"15", -- 0x0120
    x"C5",x"B8",x"A0",x"80",x"43",x"28",x"90",x"D5", -- 0x0128
    x"05",x"83",x"27",x"90",x"B8",x"3F",x"F0",x"43", -- 0x0130
    x"80",x"A0",x"14",x"E7",x"83",x"34",x"76",x"14", -- 0x0138
    x"B0",x"F2",x"3D",x"23",x"56",x"34",x"A2",x"C5", -- 0x0140
    x"FF",x"D5",x"83",x"FE",x"53",x"FE",x"AE",x"FD", -- 0x0148
    x"97",x"F7",x"F7",x"F7",x"AD",x"27",x"F7",x"4E", -- 0x0150
    x"AE",x"FC",x"67",x"37",x"17",x"6D",x"AD",x"F6", -- 0x0158
    x"6A",x"FE",x"37",x"53",x"01",x"2E",x"53",x"FE", -- 0x0160
    x"4E",x"AE",x"83",x"23",x"F8",x"B8",x"10",x"BA", -- 0x0168
    x"30",x"90",x"18",x"EA",x"71",x"83",x"A5",x"05", -- 0x0170
    x"76",x"75",x"24",x"78",x"14",x"EC",x"AA",x"B8", -- 0x0178
    x"7F",x"23",x"08",x"90",x"C8",x"F9",x"90",x"C8", -- 0x0180
    x"FA",x"47",x"53",x"0F",x"AD",x"34",x"97",x"FA", -- 0x0188
    x"53",x"0F",x"AD",x"34",x"97",x"24",x"32",x"FC", -- 0x0190
    x"90",x"C8",x"FB",x"90",x"C8",x"03",x"08",x"AB", -- 0x0198
    x"44",x"2C",x"15",x"C5",x"AC",x"BB",x"01",x"B8", -- 0x01A0
    x"3F",x"F0",x"43",x"40",x"A0",x"D5",x"05",x"83", -- 0x01A8
    x"B8",x"3E",x"F0",x"F2",x"3A",x"53",x"3F",x"D3", -- 0x01B0
    x"3B",x"96",x"3A",x"14",x"EC",x"F0",x"B8",x"02", -- 0x01B8
    x"B9",x"01",x"D2",x"E2",x"BA",x"99",x"80",x"C6", -- 0x01C0
    x"CE",x"6A",x"57",x"90",x"24",x"FC",x"81",x"C6", -- 0x01C8
    x"DA",x"23",x"59",x"90",x"81",x"6A",x"57",x"91", -- 0x01D0
    x"24",x"FC",x"B8",x"3E",x"F0",x"43",x"80",x"A0", -- 0x01D8
    x"24",x"3A",x"BA",x"01",x"80",x"D3",x"59",x"C6", -- 0x01E0
    x"EF",x"80",x"6A",x"57",x"90",x"24",x"FC",x"90", -- 0x01E8
    x"81",x"D3",x"59",x"96",x"F8",x"91",x"24",x"FC", -- 0x01F0
    x"81",x"6A",x"57",x"91",x"B8",x"7F",x"54",x"35", -- 0x01F8
    x"23",x"42",x"90",x"C8",x"B9",x"01",x"81",x"47", -- 0x0200
    x"54",x"29",x"54",x"35",x"23",x"52",x"90",x"C8", -- 0x0208
    x"81",x"54",x"29",x"54",x"35",x"23",x"56",x"90", -- 0x0210
    x"C8",x"19",x"81",x"47",x"54",x"29",x"54",x"35", -- 0x0218
    x"23",x"4A",x"90",x"C8",x"81",x"54",x"29",x"24", -- 0x0220
    x"32",x"53",x"0F",x"AD",x"34",x"4B",x"FD",x"90", -- 0x0228
    x"C8",x"FE",x"90",x"C8",x"83",x"23",x"02",x"90", -- 0x0230
    x"C8",x"83",x"B8",x"40",x"B9",x"50",x"FC",x"90", -- 0x0238
    x"91",x"18",x"19",x"FB",x"90",x"03",x"08",x"91", -- 0x0240
    x"BD",x"0A",x"B8",x"46",x"54",x"61",x"BD",x"0C", -- 0x0248
    x"B8",x"4E",x"54",x"61",x"BD",x"0C",x"B8",x"5A", -- 0x0250
    x"54",x"61",x"BD",x"0C",x"B8",x"5E",x"54",x"61", -- 0x0258
    x"83",x"34",x"4B",x"FD",x"90",x"18",x"FE",x"90", -- 0x0260
    x"18",x"83",x"07",x"BA",x"F8",x"6A",x"C9",x"F6", -- 0x0268
    x"6D",x"6A",x"53",x"07",x"17",x"AA",x"27",x"97", -- 0x0270
    x"A7",x"F7",x"EA",x"79",x"AA",x"81",x"5A",x"83", -- 0x0278
    x"54",x"6A",x"C6",x"89",x"81",x"DA",x"91",x"27", -- 0x0280
    x"17",x"83",x"54",x"6A",x"96",x"92",x"81",x"DA", -- 0x0288
    x"91",x"27",x"83",x"42",x"AC",x"53",x"0F",x"AD", -- 0x0290
    x"54",x"A4",x"2A",x"AF",x"FC",x"53",x"F0",x"47", -- 0x0298
    x"AD",x"54",x"A4",x"83",x"FD",x"03",x"B3",x"A3", -- 0x02A0
    x"96",x"AC",x"AD",x"CD",x"1D",x"AB",x"6F",x"F6", -- 0x02A8
    x"A4",x"FB",x"83",x"0F",x"0E",x"0D",x"02",x"0A", -- 0x02B0
    x"05",x"0B",x"03",x"06",x"0C",x"09",x"01",x"04", -- 0x02B8
    x"08",x"07",x"00",x"BF",x"FF",x"D5",x"14",x"F1", -- 0x02C0
    x"B9",x"F2",x"B8",x"10",x"BA",x"0B",x"BB",x"28", -- 0x02C8
    x"BC",x"70",x"BE",x"04",x"34",x"1C",x"F9",x"A3", -- 0x02D0
    x"AD",x"74",x"EA",x"19",x"1E",x"1E",x"EA",x"D6", -- 0x02D8
    x"34",x"27",x"23",x"4A",x"34",x"A2",x"34",x"3D", -- 0x02E0
    x"A9",x"34",x"1C",x"34",x"6B",x"34",x"27",x"F9", -- 0x02E8
    x"84",x"08",x"19",x"12",x"0E",x"12",x"23",x"14", -- 0x02F0
    x"0C",x"1C",x"20",x"26",x"12",x"20",x"20",x"20", -- 0x02F8
    x"00",x"0F",x"FF",x"CF",x"03",x"F0",x"3F",x"CF", -- 0x0300
    x"0F",x"0F",x"0F",x"CF",x"1C",x"71",x"C7",x"CF", -- 0x0308
    x"33",x"33",x"33",x"CF",x"03",x"F0",x"3F",x"EF", -- 0x0310
    x"0F",x"0F",x"0F",x"EF",x"1C",x"71",x"C7",x"EF", -- 0x0318
    x"33",x"33",x"33",x"EF",x"55",x"55",x"55",x"EF", -- 0x0320
    x"90",x"10",x"94",x"00",x"21",x"00",x"56",x"DF", -- 0x0328
    x"53",x"DD",x"50",x"DA",x"4D",x"D8",x"4A",x"D5", -- 0x0330
    x"47",x"D2",x"21",x"00",x"92",x"20",x"4A",x"CD", -- 0x0338
    x"52",x"EB",x"4A",x"C9",x"52",x"E7",x"4A",x"C5", -- 0x0340
    x"21",x"00",x"85",x"04",x"85",x"0C",x"85",x"14", -- 0x0348
    x"85",x"1C",x"85",x"24",x"21",x"00",x"82",x"1C", -- 0x0350
    x"21",x"00",x"8A",x"00",x"21",x"00",x"85",x"24", -- 0x0358
    x"85",x"1C",x"85",x"14",x"85",x"0C",x"85",x"04", -- 0x0360
    x"21",x"00",x"44",x"FF",x"4D",x"DD",x"48",x"DA", -- 0x0368
    x"44",x"D5",x"42",x"D3",x"21",x"00",x"F9",x"AF", -- 0x0370
    x"FE",x"39",x"FF",x"D5",x"05",x"83",x"20",x"99", -- 0x0378
    x"FE",x"84",x"08",x"99",x"FD",x"84",x"08",x"99", -- 0x0380
    x"FC",x"84",x"08",x"89",x"03",x"84",x"08",x"09", -- 0x0388
    x"A8",x"89",x"BC",x"99",x"9B",x"F9",x"43",x"F0", -- 0x0390
    x"3A",x"85",x"27",x"AA",x"AB",x"08",x"A9",x"12", -- 0x0398
    x"A2",x"CB",x"32",x"A5",x"1A",x"52",x"A8",x"1B", -- 0x03A0
    x"72",x"AB",x"CA",x"92",x"AE",x"95",x"F8",x"39", -- 0x03A8
    x"83",x"FB",x"53",x"0F",x"A8",x"FA",x"53",x"0F", -- 0x03B0
    x"47",x"48",x"A8",x"B9",x"07",x"23",x"C7",x"69", -- 0x03B8
    x"A3",x"D8",x"C6",x"C6",x"E9",x"BD",x"83",x"10", -- 0x03C0
    x"1F",x"0F",x"FF",x"F0",x"F1",x"01",x"11",x"BC", -- 0x03C8
    x"FF",x"FB",x"37",x"17",x"AE",x"FA",x"6E",x"1C", -- 0x03D0
    x"F6",x"D6",x"6B",x"AD",x"83",x"FA",x"96",x"E1", -- 0x03D8
    x"83",x"FB",x"96",x"E5",x"83",x"27",x"6B",x"EA", -- 0x03E0
    x"E6",x"83",x"FC",x"90",x"18",x"F8",x"D2",x"F9", -- 0x03E8
    x"FB",x"90",x"03",x"08",x"AB",x"18",x"54",x"61", -- 0x03F0
    x"83",x"53",x"0F",x"07",x"C6",x"F0",x"64",x"F5"  -- 0x03F8
  );

begin

  p_rom : process
  begin
    wait until rising_edge(CLK);
     D <= ROM(to_integer(unsigned(A)));
  end process;
end RTL;
