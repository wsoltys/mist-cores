-------------------------------------------------------------------------------
--
-- FPGA Videopac
--
-- $Id: mc_ctrl-c.vhd,v 1.1 2007/03/21 21:09:35 arnim Exp $
--
-------------------------------------------------------------------------------

configuration mc_ctrl_rtl_c0 of mc_ctrl is

  for rtl
  end for;

end mc_ctrl_rtl_c0;
