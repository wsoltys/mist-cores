-------------------------------------------------------------------------------
--
-- FPGA Videopac
--
-- $Id: dpram-c.vhd,v 1.1 2007/01/05 21:55:11 arnim Exp $
--
-------------------------------------------------------------------------------

configuration dpram_rtl_c0 of dpram is

  for rtl
  end for;

end dpram_rtl_c0;
