-------------------------------------------------------------------------------
--
-- FPGA Videopac
--
-- $Id: vp_por-c.vhd,v 1.2 2007/01/05 22:02:59 arnim Exp $
--
-------------------------------------------------------------------------------

configuration vp_por_rtl_c0 of vp_por is

  for spartan
  end for;

end vp_por_rtl_c0;
